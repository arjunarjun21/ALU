* NGSPICE file created from alu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

.subckt alu A[0] A[1] A[2] A[3] B[0] B[1] B[2] B[3] SEL[0] SEL[1] VGND VPWR Y[0] Y[1]
+ Y[2] Y[3]
XTAP_TAPCELL_ROW_8_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_49_ net3 _16_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_48_ net7 _15_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 net6 _05_ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput11 net11 VGND VGND VPWR VPWR Y[0] sky130_fd_sc_hd__buf_2
X_63_ _01_ _21_ _28_ net10 _29_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__o221a_1
X_46_ _04_ _09_ _08_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput12 net12 VGND VGND VPWR VPWR Y[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_62_ net10 _24_ VGND VGND VPWR VPWR _29_ sky130_fd_sc_hd__nand2_1
X_45_ net6 _01_ _12_ _13_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__o211a_1
Xoutput13 net13 VGND VGND VPWR VPWR Y[2] sky130_fd_sc_hd__clkbuf_4
X_61_ _23_ _27_ VGND VGND VPWR VPWR _28_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_44_ net9 net6 net2 _00_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput14 net14 VGND VGND VPWR VPWR Y[3] sky130_fd_sc_hd__buf_2
X_60_ _25_ _26_ VGND VGND VPWR VPWR _27_ sky130_fd_sc_hd__xnor2_1
X_43_ _00_ _11_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_42_ _04_ _10_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_41_ _08_ _09_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_40_ net2 _06_ _07_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 A[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 A[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_0_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 A[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 A[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 B[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_3_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_59_ net5 net6 net7 _05_ VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 B[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
X_58_ _24_ _21_ VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 B[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_57_ net8 net4 VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__nor2_1
Xinput10 SEL[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_56_ _14_ _17_ _22_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__a21oi_1
Xinput8 B[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_39_ _06_ _07_ net2 VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 SEL[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_0_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ _16_ net3 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__and2b_1
X_38_ net5 _05_ net6 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_54_ net8 net4 VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_37_ net5 net6 _05_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_53_ net3 _01_ _19_ _20_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_7_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36_ net10 net9 VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_52_ net9 net3 net7 _00_ VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__a211o_1
X_35_ net1 net5 VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_51_ _00_ _18_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__nand2_1
X_34_ net1 net5 _03_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__o21a_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_50_ _14_ _17_ VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__xnor2_1
X_33_ net10 _01_ _02_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net1 net5 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31_ _00_ net9 VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30_ net10 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

