VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu
  CLASS BLOCK ;
  FOREIGN alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 44.095 BY 54.815 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 40.095 13.640 44.095 14.240 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 40.095 30.640 44.095 31.240 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END A[3]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 40.095 23.840 44.095 24.440 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 40.095 37.440 44.095 38.040 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END B[3]
  PIN SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 40.095 27.240 44.095 27.840 ;
    END
  END SEL[0]
  PIN SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 40.095 20.440 44.095 21.040 ;
    END
  END SEL[1]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.100 10.640 13.700 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.265 10.640 21.865 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.430 10.640 30.030 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.595 10.640 38.195 43.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.460 38.420 19.060 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 25.620 38.420 27.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 33.780 38.420 35.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.940 38.420 43.540 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.800 10.640 10.400 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.965 10.640 18.565 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.130 10.640 26.730 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.295 10.640 34.895 43.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.160 38.420 15.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 22.320 38.420 23.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.480 38.420 32.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 38.640 38.420 40.240 ;
    END
  END VPWR
  PIN Y[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 40.095 17.040 44.095 17.640 ;
    END
  END Y[0]
  PIN Y[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 40.095 34.040 44.095 34.640 ;
    END
  END Y[1]
  PIN Y[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 50.815 19.690 54.815 ;
    END
  END Y[2]
  PIN Y[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END Y[3]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 38.370 43.605 ;
      LAYER li1 ;
        RECT 5.520 10.795 38.180 43.605 ;
      LAYER met1 ;
        RECT 4.210 10.640 39.030 43.760 ;
      LAYER met2 ;
        RECT 4.230 50.535 19.130 51.410 ;
        RECT 19.970 50.535 39.010 51.410 ;
        RECT 4.230 4.280 39.010 50.535 ;
        RECT 4.230 3.670 12.690 4.280 ;
        RECT 13.530 3.670 15.910 4.280 ;
        RECT 16.750 3.670 19.130 4.280 ;
        RECT 19.970 3.670 39.010 4.280 ;
      LAYER met3 ;
        RECT 3.990 38.440 40.095 43.685 ;
        RECT 3.990 37.040 39.695 38.440 ;
        RECT 3.990 35.040 40.095 37.040 ;
        RECT 4.400 33.640 39.695 35.040 ;
        RECT 3.990 31.640 40.095 33.640 ;
        RECT 4.400 30.240 39.695 31.640 ;
        RECT 3.990 28.240 40.095 30.240 ;
        RECT 3.990 26.840 39.695 28.240 ;
        RECT 3.990 24.840 40.095 26.840 ;
        RECT 3.990 23.440 39.695 24.840 ;
        RECT 3.990 21.440 40.095 23.440 ;
        RECT 3.990 20.040 39.695 21.440 ;
        RECT 3.990 18.040 40.095 20.040 ;
        RECT 3.990 16.640 39.695 18.040 ;
        RECT 3.990 14.640 40.095 16.640 ;
        RECT 3.990 13.240 39.695 14.640 ;
        RECT 3.990 10.715 40.095 13.240 ;
  END
END alu
END LIBRARY

