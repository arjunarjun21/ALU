magic
tech sky130A
magscale 1 2
timestamp 1752153290
<< checkpaint >>
rect -3932 -3932 12751 14895
<< viali >>
rect 3985 8517 4019 8551
rect 4353 8449 4387 8483
rect 7021 7837 7055 7871
rect 7297 7837 7331 7871
rect 1409 7361 1443 7395
rect 2513 7361 2547 7395
rect 3341 7361 3375 7395
rect 3525 7361 3559 7395
rect 5733 7361 5767 7395
rect 7021 7361 7055 7395
rect 2605 7293 2639 7327
rect 5825 7293 5859 7327
rect 2881 7225 2915 7259
rect 6101 7225 6135 7259
rect 1593 7157 1627 7191
rect 3433 7157 3467 7191
rect 7205 7157 7239 7191
rect 6101 6953 6135 6987
rect 3065 6885 3099 6919
rect 3249 6885 3283 6919
rect 6285 6885 6319 6919
rect 2145 6817 2179 6851
rect 4445 6817 4479 6851
rect 6009 6817 6043 6851
rect 2237 6749 2271 6783
rect 3525 6749 3559 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4997 6749 5031 6783
rect 5273 6749 5307 6783
rect 5365 6749 5399 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 5733 6749 5767 6783
rect 6653 6749 6687 6783
rect 6837 6749 6871 6783
rect 2697 6681 2731 6715
rect 3249 6681 3283 6715
rect 3433 6681 3467 6715
rect 6561 6681 6595 6715
rect 2605 6613 2639 6647
rect 3157 6613 3191 6647
rect 4813 6613 4847 6647
rect 5181 6613 5215 6647
rect 6653 6613 6687 6647
rect 3801 6409 3835 6443
rect 4997 6409 5031 6443
rect 5641 6409 5675 6443
rect 6745 6409 6779 6443
rect 4905 6341 4939 6375
rect 1409 6273 1443 6307
rect 3249 6273 3283 6307
rect 3341 6273 3375 6307
rect 3525 6273 3559 6307
rect 3617 6273 3651 6307
rect 4721 6273 4755 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 7297 6273 7331 6307
rect 6101 6205 6135 6239
rect 6469 6205 6503 6239
rect 1593 6137 1627 6171
rect 7113 6137 7147 6171
rect 4537 6069 4571 6103
rect 6009 6069 6043 6103
rect 6377 6069 6411 6103
rect 2329 5865 2363 5899
rect 7113 5797 7147 5831
rect 2697 5729 2731 5763
rect 2605 5661 2639 5695
rect 7297 5661 7331 5695
rect 4261 5321 4295 5355
rect 4813 5321 4847 5355
rect 5825 5321 5859 5355
rect 5457 5253 5491 5287
rect 5657 5253 5691 5287
rect 6009 5253 6043 5287
rect 7021 5253 7055 5287
rect 4537 5185 4571 5219
rect 4905 5185 4939 5219
rect 5917 5185 5951 5219
rect 6193 5185 6227 5219
rect 7205 5185 7239 5219
rect 4261 5117 4295 5151
rect 4445 5049 4479 5083
rect 6193 5049 6227 5083
rect 5641 4981 5675 5015
rect 4813 4777 4847 4811
rect 5181 4777 5215 4811
rect 4169 4709 4203 4743
rect 4261 4709 4295 4743
rect 7021 4641 7055 4675
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 5273 4573 5307 4607
rect 7297 4573 7331 4607
rect 3893 4437 3927 4471
rect 2697 4097 2731 4131
rect 2881 4097 2915 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 2881 3893 2915 3927
rect 5733 3893 5767 3927
rect 6009 3689 6043 3723
rect 6193 3689 6227 3723
rect 3065 3621 3099 3655
rect 2697 3553 2731 3587
rect 3525 3553 3559 3587
rect 4169 3553 4203 3587
rect 5733 3553 5767 3587
rect 2145 3485 2179 3519
rect 2329 3485 2363 3519
rect 2605 3485 2639 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4353 3485 4387 3519
rect 5641 3485 5675 3519
rect 6469 3485 6503 3519
rect 7021 3485 7055 3519
rect 5549 3417 5583 3451
rect 2237 3349 2271 3383
rect 2973 3349 3007 3383
rect 4537 3349 4571 3383
rect 5181 3349 5215 3383
rect 7205 3349 7239 3383
rect 2973 3145 3007 3179
rect 3249 3145 3283 3179
rect 5273 3145 5307 3179
rect 2605 3009 2639 3043
rect 2789 3009 2823 3043
rect 3065 3009 3099 3043
rect 3249 3009 3283 3043
rect 5457 3009 5491 3043
rect 5641 3009 5675 3043
rect 7297 3009 7331 3043
rect 5733 2941 5767 2975
rect 7113 2873 7147 2907
rect 2697 2601 2731 2635
rect 3341 2601 3375 2635
rect 2881 2397 2915 2431
rect 3525 2397 3559 2431
rect 4261 2397 4295 2431
rect 4077 2261 4111 2295
<< metal1 >>
rect 1104 8730 7639 8752
rect 1104 8678 2426 8730
rect 2478 8678 2490 8730
rect 2542 8678 2554 8730
rect 2606 8678 2618 8730
rect 2670 8678 2682 8730
rect 2734 8678 4059 8730
rect 4111 8678 4123 8730
rect 4175 8678 4187 8730
rect 4239 8678 4251 8730
rect 4303 8678 4315 8730
rect 4367 8678 5692 8730
rect 5744 8678 5756 8730
rect 5808 8678 5820 8730
rect 5872 8678 5884 8730
rect 5936 8678 5948 8730
rect 6000 8678 7325 8730
rect 7377 8678 7389 8730
rect 7441 8678 7453 8730
rect 7505 8678 7517 8730
rect 7569 8678 7581 8730
rect 7633 8678 7639 8730
rect 1104 8656 7639 8678
rect 3970 8508 3976 8560
rect 4028 8508 4034 8560
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4430 8480 4436 8492
rect 4387 8452 4436 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 1104 8186 7636 8208
rect 1104 8134 1766 8186
rect 1818 8134 1830 8186
rect 1882 8134 1894 8186
rect 1946 8134 1958 8186
rect 2010 8134 2022 8186
rect 2074 8134 3399 8186
rect 3451 8134 3463 8186
rect 3515 8134 3527 8186
rect 3579 8134 3591 8186
rect 3643 8134 3655 8186
rect 3707 8134 5032 8186
rect 5084 8134 5096 8186
rect 5148 8134 5160 8186
rect 5212 8134 5224 8186
rect 5276 8134 5288 8186
rect 5340 8134 6665 8186
rect 6717 8134 6729 8186
rect 6781 8134 6793 8186
rect 6845 8134 6857 8186
rect 6909 8134 6921 8186
rect 6973 8134 7636 8186
rect 1104 8112 7636 8134
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6236 7840 7021 7868
rect 6236 7828 6242 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 7742 7868 7748 7880
rect 7331 7840 7748 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 1104 7642 7639 7664
rect 1104 7590 2426 7642
rect 2478 7590 2490 7642
rect 2542 7590 2554 7642
rect 2606 7590 2618 7642
rect 2670 7590 2682 7642
rect 2734 7590 4059 7642
rect 4111 7590 4123 7642
rect 4175 7590 4187 7642
rect 4239 7590 4251 7642
rect 4303 7590 4315 7642
rect 4367 7590 5692 7642
rect 5744 7590 5756 7642
rect 5808 7590 5820 7642
rect 5872 7590 5884 7642
rect 5936 7590 5948 7642
rect 6000 7590 7325 7642
rect 7377 7590 7389 7642
rect 7441 7590 7453 7642
rect 7505 7590 7517 7642
rect 7569 7590 7581 7642
rect 7633 7590 7639 7642
rect 1104 7568 7639 7590
rect 3234 7460 3240 7472
rect 2746 7432 3240 7460
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2746 7392 2774 7432
rect 3234 7420 3240 7432
rect 3292 7420 3298 7472
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 2547 7364 2774 7392
rect 2884 7364 3341 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2590 7284 2596 7336
rect 2648 7284 2654 7336
rect 2884 7265 2912 7364
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3878 7392 3884 7404
rect 3559 7364 3884 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5592 7364 5733 7392
rect 5592 7352 5598 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6052 7364 7021 7392
rect 6052 7352 6058 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 5810 7284 5816 7336
rect 5868 7284 5874 7336
rect 2869 7259 2927 7265
rect 2869 7225 2881 7259
rect 2915 7225 2927 7259
rect 2869 7219 2927 7225
rect 6086 7216 6092 7268
rect 6144 7216 6150 7268
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 2222 7188 2228 7200
rect 1627 7160 2228 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 3970 7188 3976 7200
rect 3467 7160 3976 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 6178 7188 6184 7200
rect 5776 7160 6184 7188
rect 5776 7148 5782 7160
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 7190 7148 7196 7200
rect 7248 7148 7254 7200
rect 1104 7098 7636 7120
rect 1104 7046 1766 7098
rect 1818 7046 1830 7098
rect 1882 7046 1894 7098
rect 1946 7046 1958 7098
rect 2010 7046 2022 7098
rect 2074 7046 3399 7098
rect 3451 7046 3463 7098
rect 3515 7046 3527 7098
rect 3579 7046 3591 7098
rect 3643 7046 3655 7098
rect 3707 7046 5032 7098
rect 5084 7046 5096 7098
rect 5148 7046 5160 7098
rect 5212 7046 5224 7098
rect 5276 7046 5288 7098
rect 5340 7046 6665 7098
rect 6717 7046 6729 7098
rect 6781 7046 6793 7098
rect 6845 7046 6857 7098
rect 6909 7046 6921 7098
rect 6973 7046 7636 7098
rect 1104 7024 7636 7046
rect 3068 6956 3372 6984
rect 3068 6925 3096 6956
rect 3053 6919 3111 6925
rect 3053 6885 3065 6919
rect 3099 6885 3111 6919
rect 3053 6879 3111 6885
rect 3237 6919 3295 6925
rect 3237 6885 3249 6919
rect 3283 6885 3295 6919
rect 3237 6879 3295 6885
rect 2130 6808 2136 6860
rect 2188 6808 2194 6860
rect 3068 6848 3096 6879
rect 2240 6820 3096 6848
rect 2240 6792 2268 6820
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 3252 6848 3280 6879
rect 3200 6820 3280 6848
rect 3344 6848 3372 6956
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 5868 6956 6101 6984
rect 5868 6944 5874 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 6273 6919 6331 6925
rect 6273 6916 6285 6919
rect 5316 6888 6285 6916
rect 5316 6876 5322 6888
rect 6273 6885 6285 6888
rect 6319 6916 6331 6919
rect 6638 6916 6644 6928
rect 6319 6888 6644 6916
rect 6319 6885 6331 6888
rect 6273 6879 6331 6885
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 3344 6820 3648 6848
rect 3200 6808 3206 6820
rect 2222 6740 2228 6792
rect 2280 6740 2286 6792
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 2648 6752 3525 6780
rect 2648 6740 2654 6752
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3620 6724 3648 6820
rect 4080 6820 4292 6848
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4080 6789 4108 6820
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4264 6780 4292 6820
rect 4430 6808 4436 6860
rect 4488 6808 4494 6860
rect 5000 6820 5856 6848
rect 4614 6780 4620 6792
rect 4264 6752 4620 6780
rect 4157 6743 4215 6749
rect 2130 6672 2136 6724
rect 2188 6712 2194 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2188 6684 2697 6712
rect 2188 6672 2194 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 3237 6715 3295 6721
rect 3237 6681 3249 6715
rect 3283 6681 3295 6715
rect 3237 6675 3295 6681
rect 2590 6604 2596 6656
rect 2648 6604 2654 6656
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3252 6644 3280 6675
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 3421 6715 3479 6721
rect 3421 6712 3433 6715
rect 3384 6684 3433 6712
rect 3384 6672 3390 6684
rect 3421 6681 3433 6684
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 3191 6616 3280 6644
rect 3436 6644 3464 6675
rect 3602 6672 3608 6724
rect 3660 6712 3666 6724
rect 4172 6712 4200 6743
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5000 6789 5028 6820
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 5460 6752 5549 6780
rect 3660 6684 4200 6712
rect 5460 6712 5488 6752
rect 5537 6749 5549 6752
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5828 6780 5856 6820
rect 5994 6808 6000 6860
rect 6052 6808 6058 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6144 6820 6868 6848
rect 6144 6808 6150 6820
rect 6641 6783 6699 6789
rect 5828 6752 6592 6780
rect 6564 6724 6592 6752
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 6730 6780 6736 6792
rect 6687 6752 6736 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 6840 6789 6868 6820
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 5460 6684 5575 6712
rect 3660 6672 3666 6684
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 3436 6616 4813 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5442 6644 5448 6656
rect 5215 6616 5448 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5547 6644 5575 6684
rect 6546 6672 6552 6724
rect 6604 6672 6610 6724
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 5547 6616 6653 6644
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6641 6607 6699 6613
rect 1104 6554 7639 6576
rect 1104 6502 2426 6554
rect 2478 6502 2490 6554
rect 2542 6502 2554 6554
rect 2606 6502 2618 6554
rect 2670 6502 2682 6554
rect 2734 6502 4059 6554
rect 4111 6502 4123 6554
rect 4175 6502 4187 6554
rect 4239 6502 4251 6554
rect 4303 6502 4315 6554
rect 4367 6502 5692 6554
rect 5744 6502 5756 6554
rect 5808 6502 5820 6554
rect 5872 6502 5884 6554
rect 5936 6502 5948 6554
rect 6000 6502 7325 6554
rect 7377 6502 7389 6554
rect 7441 6502 7453 6554
rect 7505 6502 7517 6554
rect 7569 6502 7581 6554
rect 7633 6502 7639 6554
rect 1104 6480 7639 6502
rect 3786 6400 3792 6452
rect 3844 6400 3850 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5350 6440 5356 6452
rect 5031 6412 5356 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 6546 6440 6552 6452
rect 5675 6412 6552 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6696 6412 6745 6440
rect 6696 6400 6702 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 4893 6375 4951 6381
rect 4893 6372 4905 6375
rect 3528 6344 4905 6372
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 3234 6264 3240 6316
rect 3292 6264 3298 6316
rect 3528 6313 3556 6344
rect 4893 6341 4905 6344
rect 4939 6372 4951 6375
rect 4939 6344 5304 6372
rect 4939 6341 4951 6344
rect 4893 6335 4951 6341
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3344 6236 3372 6267
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 5276 6313 5304 6344
rect 5460 6344 6500 6372
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5350 6304 5356 6316
rect 5307 6276 5356 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 4522 6236 4528 6248
rect 1596 6208 4528 6236
rect 1596 6177 1624 6208
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6137 1639 6171
rect 1581 6131 1639 6137
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 3878 6168 3884 6180
rect 3292 6140 3884 6168
rect 3292 6128 3298 6140
rect 3878 6128 3884 6140
rect 3936 6168 3942 6180
rect 4724 6168 4752 6267
rect 5184 6236 5212 6267
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5460 6313 5488 6344
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5718 6304 5724 6316
rect 5583 6276 5724 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5828 6313 5856 6344
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6236 6276 6377 6304
rect 6236 6264 6242 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 5994 6236 6000 6248
rect 5184 6208 6000 6236
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6086 6196 6092 6248
rect 6144 6196 6150 6248
rect 6472 6245 6500 6344
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6236 6515 6239
rect 6503 6208 7144 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 4798 6168 4804 6180
rect 3936 6140 4804 6168
rect 3936 6128 3942 6140
rect 4798 6128 4804 6140
rect 4856 6168 4862 6180
rect 5718 6168 5724 6180
rect 4856 6140 5724 6168
rect 4856 6128 4862 6140
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 6104 6168 6132 6196
rect 7116 6177 7144 6208
rect 7101 6171 7159 6177
rect 6104 6140 6408 6168
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4614 6100 4620 6112
rect 4571 6072 4620 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5997 6103 6055 6109
rect 5997 6069 6009 6103
rect 6043 6100 6055 6103
rect 6178 6100 6184 6112
rect 6043 6072 6184 6100
rect 6043 6069 6055 6072
rect 5997 6063 6055 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6380 6109 6408 6140
rect 7101 6137 7113 6171
rect 7147 6137 7159 6171
rect 7101 6131 7159 6137
rect 6365 6103 6423 6109
rect 6365 6069 6377 6103
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 1104 6010 7636 6032
rect 1104 5958 1766 6010
rect 1818 5958 1830 6010
rect 1882 5958 1894 6010
rect 1946 5958 1958 6010
rect 2010 5958 2022 6010
rect 2074 5958 3399 6010
rect 3451 5958 3463 6010
rect 3515 5958 3527 6010
rect 3579 5958 3591 6010
rect 3643 5958 3655 6010
rect 3707 5958 5032 6010
rect 5084 5958 5096 6010
rect 5148 5958 5160 6010
rect 5212 5958 5224 6010
rect 5276 5958 5288 6010
rect 5340 5958 6665 6010
rect 6717 5958 6729 6010
rect 6781 5958 6793 6010
rect 6845 5958 6857 6010
rect 6909 5958 6921 6010
rect 6973 5958 7636 6010
rect 1104 5936 7636 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 2188 5868 2329 5896
rect 2188 5856 2194 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 2317 5859 2375 5865
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 7101 5831 7159 5837
rect 7101 5828 7113 5831
rect 5408 5800 7113 5828
rect 5408 5788 5414 5800
rect 7101 5797 7113 5800
rect 7147 5797 7159 5831
rect 7101 5791 7159 5797
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 4430 5760 4436 5772
rect 2731 5732 4436 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 4522 5692 4528 5704
rect 2639 5664 4528 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7742 5692 7748 5704
rect 7331 5664 7748 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 1104 5466 7639 5488
rect 1104 5414 2426 5466
rect 2478 5414 2490 5466
rect 2542 5414 2554 5466
rect 2606 5414 2618 5466
rect 2670 5414 2682 5466
rect 2734 5414 4059 5466
rect 4111 5414 4123 5466
rect 4175 5414 4187 5466
rect 4239 5414 4251 5466
rect 4303 5414 4315 5466
rect 4367 5414 5692 5466
rect 5744 5414 5756 5466
rect 5808 5414 5820 5466
rect 5872 5414 5884 5466
rect 5936 5414 5948 5466
rect 6000 5414 7325 5466
rect 7377 5414 7389 5466
rect 7441 5414 7453 5466
rect 7505 5414 7517 5466
rect 7569 5414 7581 5466
rect 7633 5414 7639 5466
rect 1104 5392 7639 5414
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4430 5352 4436 5364
rect 4295 5324 4436 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 4798 5312 4804 5364
rect 4856 5312 4862 5364
rect 5813 5355 5871 5361
rect 5460 5324 5764 5352
rect 5460 5293 5488 5324
rect 5445 5287 5503 5293
rect 5445 5284 5457 5287
rect 4540 5256 5457 5284
rect 4540 5225 4568 5256
rect 5445 5253 5457 5256
rect 5491 5253 5503 5287
rect 5645 5287 5703 5293
rect 5645 5284 5657 5287
rect 5445 5247 5503 5253
rect 5644 5253 5657 5284
rect 5691 5253 5703 5287
rect 5736 5284 5764 5324
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 6086 5352 6092 5364
rect 5859 5324 6092 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 5997 5287 6055 5293
rect 5997 5284 6009 5287
rect 5736 5256 6009 5284
rect 5644 5247 5703 5253
rect 5997 5253 6009 5256
rect 6043 5284 6055 5287
rect 7009 5287 7067 5293
rect 7009 5284 7021 5287
rect 6043 5256 7021 5284
rect 6043 5253 6055 5256
rect 5997 5247 6055 5253
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4798 5148 4804 5160
rect 4295 5120 4804 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4798 5108 4804 5120
rect 4856 5148 4862 5160
rect 5644 5148 5672 5247
rect 6104 5228 6132 5256
rect 7009 5253 7021 5256
rect 7055 5253 7067 5287
rect 7009 5247 7067 5253
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 5920 5148 5948 5179
rect 6086 5176 6092 5228
rect 6144 5176 6150 5228
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6270 5216 6276 5228
rect 6227 5188 6276 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 7190 5176 7196 5228
rect 7248 5176 7254 5228
rect 4856 5120 5948 5148
rect 4856 5108 4862 5120
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4433 5083 4491 5089
rect 4433 5080 4445 5083
rect 4212 5052 4445 5080
rect 4212 5040 4218 5052
rect 4433 5049 4445 5052
rect 4479 5080 4491 5083
rect 4479 5052 5672 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 5644 5021 5672 5052
rect 6178 5040 6184 5092
rect 6236 5040 6242 5092
rect 5629 5015 5687 5021
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 6270 5012 6276 5024
rect 5675 4984 6276 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 1104 4922 7636 4944
rect 1104 4870 1766 4922
rect 1818 4870 1830 4922
rect 1882 4870 1894 4922
rect 1946 4870 1958 4922
rect 2010 4870 2022 4922
rect 2074 4870 3399 4922
rect 3451 4870 3463 4922
rect 3515 4870 3527 4922
rect 3579 4870 3591 4922
rect 3643 4870 3655 4922
rect 3707 4870 5032 4922
rect 5084 4870 5096 4922
rect 5148 4870 5160 4922
rect 5212 4870 5224 4922
rect 5276 4870 5288 4922
rect 5340 4870 6665 4922
rect 6717 4870 6729 4922
rect 6781 4870 6793 4922
rect 6845 4870 6857 4922
rect 6909 4870 6921 4922
rect 6973 4870 7636 4922
rect 1104 4848 7636 4870
rect 4798 4768 4804 4820
rect 4856 4768 4862 4820
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4948 4780 5181 4808
rect 4948 4768 4954 4780
rect 5169 4777 5181 4780
rect 5215 4808 5227 4811
rect 5350 4808 5356 4820
rect 5215 4780 5356 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5350 4768 5356 4780
rect 5408 4808 5414 4820
rect 5408 4780 7052 4808
rect 5408 4768 5414 4780
rect 4154 4700 4160 4752
rect 4212 4700 4218 4752
rect 4249 4743 4307 4749
rect 4249 4709 4261 4743
rect 4295 4740 4307 4743
rect 4522 4740 4528 4752
rect 4295 4712 4528 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 4816 4672 4844 4768
rect 7024 4681 7052 4780
rect 4356 4644 4844 4672
rect 7009 4675 7067 4681
rect 4356 4613 4384 4644
rect 7009 4641 7021 4675
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5442 4604 5448 4616
rect 5307 4576 5448 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 4080 4536 4108 4567
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7742 4604 7748 4616
rect 7331 4576 7748 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 6086 4536 6092 4548
rect 4080 4508 6092 4536
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 3878 4428 3884 4480
rect 3936 4428 3942 4480
rect 1104 4378 7639 4400
rect 1104 4326 2426 4378
rect 2478 4326 2490 4378
rect 2542 4326 2554 4378
rect 2606 4326 2618 4378
rect 2670 4326 2682 4378
rect 2734 4326 4059 4378
rect 4111 4326 4123 4378
rect 4175 4326 4187 4378
rect 4239 4326 4251 4378
rect 4303 4326 4315 4378
rect 4367 4326 5692 4378
rect 5744 4326 5756 4378
rect 5808 4326 5820 4378
rect 5872 4326 5884 4378
rect 5936 4326 5948 4378
rect 6000 4326 7325 4378
rect 7377 4326 7389 4378
rect 7441 4326 7453 4378
rect 7505 4326 7517 4378
rect 7569 4326 7581 4378
rect 7633 4326 7639 4378
rect 1104 4304 7639 4326
rect 6086 4196 6092 4208
rect 5644 4168 6092 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2774 4128 2780 4140
rect 2731 4100 2780 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 2958 4128 2964 4140
rect 2915 4100 2964 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 5644 4137 5672 4168
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6178 4128 6184 4140
rect 5859 4100 6184 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 5718 3884 5724 3936
rect 5776 3884 5782 3936
rect 1104 3834 7636 3856
rect 1104 3782 1766 3834
rect 1818 3782 1830 3834
rect 1882 3782 1894 3834
rect 1946 3782 1958 3834
rect 2010 3782 2022 3834
rect 2074 3782 3399 3834
rect 3451 3782 3463 3834
rect 3515 3782 3527 3834
rect 3579 3782 3591 3834
rect 3643 3782 3655 3834
rect 3707 3782 5032 3834
rect 5084 3782 5096 3834
rect 5148 3782 5160 3834
rect 5212 3782 5224 3834
rect 5276 3782 5288 3834
rect 5340 3782 6665 3834
rect 6717 3782 6729 3834
rect 6781 3782 6793 3834
rect 6845 3782 6857 3834
rect 6909 3782 6921 3834
rect 6973 3782 7636 3834
rect 1104 3760 7636 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3016 3692 4016 3720
rect 3016 3680 3022 3692
rect 3053 3655 3111 3661
rect 3053 3652 3065 3655
rect 2700 3624 3065 3652
rect 2700 3593 2728 3624
rect 3053 3621 3065 3624
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3553 2743 3587
rect 3142 3584 3148 3596
rect 2685 3547 2743 3553
rect 2792 3556 3148 3584
rect 2130 3476 2136 3528
rect 2188 3476 2194 3528
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2792 3516 2820 3556
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 3878 3584 3884 3596
rect 3559 3556 3884 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 3988 3584 4016 3692
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5592 3692 6009 3720
rect 5592 3680 5598 3692
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 5997 3683 6055 3689
rect 6178 3680 6184 3732
rect 6236 3680 6242 3732
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 3988 3556 4169 3584
rect 4157 3553 4169 3556
rect 4203 3553 4215 3587
rect 4157 3547 4215 3553
rect 5718 3544 5724 3596
rect 5776 3544 5782 3596
rect 2639 3488 2820 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 2924 3488 3433 3516
rect 2924 3476 2930 3488
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4614 3516 4620 3528
rect 4387 3488 4620 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 3988 3448 4016 3479
rect 2976 3420 4016 3448
rect 4080 3448 4108 3479
rect 4614 3476 4620 3488
rect 4672 3516 4678 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 4672 3488 5641 3516
rect 4672 3476 4678 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6144 3488 6469 3516
rect 6144 3476 6150 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 7006 3476 7012 3528
rect 7064 3476 7070 3528
rect 4430 3448 4436 3460
rect 4080 3420 4436 3448
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3380 2283 3383
rect 2866 3380 2872 3392
rect 2271 3352 2872 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 2976 3389 3004 3420
rect 4430 3408 4436 3420
rect 4488 3448 4494 3460
rect 5350 3448 5356 3460
rect 4488 3420 5356 3448
rect 4488 3408 4494 3420
rect 5350 3408 5356 3420
rect 5408 3448 5414 3460
rect 5537 3451 5595 3457
rect 5537 3448 5549 3451
rect 5408 3420 5549 3448
rect 5408 3408 5414 3420
rect 5537 3417 5549 3420
rect 5583 3417 5595 3451
rect 5537 3411 5595 3417
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 5169 3383 5227 3389
rect 5169 3349 5181 3383
rect 5215 3380 5227 3383
rect 5442 3380 5448 3392
rect 5215 3352 5448 3380
rect 5215 3349 5227 3352
rect 5169 3343 5227 3349
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 1104 3290 7639 3312
rect 1104 3238 2426 3290
rect 2478 3238 2490 3290
rect 2542 3238 2554 3290
rect 2606 3238 2618 3290
rect 2670 3238 2682 3290
rect 2734 3238 4059 3290
rect 4111 3238 4123 3290
rect 4175 3238 4187 3290
rect 4239 3238 4251 3290
rect 4303 3238 4315 3290
rect 4367 3238 5692 3290
rect 5744 3238 5756 3290
rect 5808 3238 5820 3290
rect 5872 3238 5884 3290
rect 5936 3238 5948 3290
rect 6000 3238 7325 3290
rect 7377 3238 7389 3290
rect 7441 3238 7453 3290
rect 7505 3238 7517 3290
rect 7569 3238 7581 3290
rect 7633 3238 7639 3290
rect 1104 3216 7639 3238
rect 2774 3176 2780 3188
rect 2746 3136 2780 3176
rect 2832 3136 2838 3188
rect 2958 3136 2964 3188
rect 3016 3136 3022 3188
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 3786 3176 3792 3188
rect 3283 3148 3792 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 7006 3176 7012 3188
rect 5307 3148 7012 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 2314 3068 2320 3120
rect 2372 3108 2378 3120
rect 2746 3108 2774 3136
rect 2372 3080 2774 3108
rect 2372 3068 2378 3080
rect 2866 3068 2872 3120
rect 2924 3108 2930 3120
rect 2924 3080 3096 3108
rect 2924 3068 2930 3080
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2188 3012 2605 3040
rect 2188 3000 2194 3012
rect 2593 3009 2605 3012
rect 2639 3040 2651 3043
rect 2682 3040 2688 3052
rect 2639 3012 2688 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 3068 3049 3096 3080
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 4430 3040 4436 3052
rect 3283 3012 4436 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 6086 3040 6092 3052
rect 5675 3012 6092 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 7282 3000 7288 3052
rect 7340 3000 7346 3052
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2941 5779 2975
rect 5721 2935 5779 2941
rect 5736 2904 5764 2935
rect 6178 2904 6184 2916
rect 5736 2876 6184 2904
rect 6178 2864 6184 2876
rect 6236 2904 6242 2916
rect 7101 2907 7159 2913
rect 7101 2904 7113 2907
rect 6236 2876 7113 2904
rect 6236 2864 6242 2876
rect 7101 2873 7113 2876
rect 7147 2873 7159 2907
rect 7101 2867 7159 2873
rect 1104 2746 7636 2768
rect 1104 2694 1766 2746
rect 1818 2694 1830 2746
rect 1882 2694 1894 2746
rect 1946 2694 1958 2746
rect 2010 2694 2022 2746
rect 2074 2694 3399 2746
rect 3451 2694 3463 2746
rect 3515 2694 3527 2746
rect 3579 2694 3591 2746
rect 3643 2694 3655 2746
rect 3707 2694 5032 2746
rect 5084 2694 5096 2746
rect 5148 2694 5160 2746
rect 5212 2694 5224 2746
rect 5276 2694 5288 2746
rect 5340 2694 6665 2746
rect 6717 2694 6729 2746
rect 6781 2694 6793 2746
rect 6845 2694 6857 2746
rect 6909 2694 6921 2746
rect 6973 2694 7636 2746
rect 1104 2672 7636 2694
rect 2682 2592 2688 2644
rect 2740 2592 2746 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 2832 2604 3341 2632
rect 2832 2592 2838 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 3329 2595 3387 2601
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2372 2400 2881 2428
rect 2372 2388 2378 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3292 2400 3525 2428
rect 3292 2388 3298 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4522 2428 4528 2440
rect 4295 2400 4528 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 1104 2202 7639 2224
rect 1104 2150 2426 2202
rect 2478 2150 2490 2202
rect 2542 2150 2554 2202
rect 2606 2150 2618 2202
rect 2670 2150 2682 2202
rect 2734 2150 4059 2202
rect 4111 2150 4123 2202
rect 4175 2150 4187 2202
rect 4239 2150 4251 2202
rect 4303 2150 4315 2202
rect 4367 2150 5692 2202
rect 5744 2150 5756 2202
rect 5808 2150 5820 2202
rect 5872 2150 5884 2202
rect 5936 2150 5948 2202
rect 6000 2150 7325 2202
rect 7377 2150 7389 2202
rect 7441 2150 7453 2202
rect 7505 2150 7517 2202
rect 7569 2150 7581 2202
rect 7633 2150 7639 2202
rect 1104 2128 7639 2150
<< via1 >>
rect 2426 8678 2478 8730
rect 2490 8678 2542 8730
rect 2554 8678 2606 8730
rect 2618 8678 2670 8730
rect 2682 8678 2734 8730
rect 4059 8678 4111 8730
rect 4123 8678 4175 8730
rect 4187 8678 4239 8730
rect 4251 8678 4303 8730
rect 4315 8678 4367 8730
rect 5692 8678 5744 8730
rect 5756 8678 5808 8730
rect 5820 8678 5872 8730
rect 5884 8678 5936 8730
rect 5948 8678 6000 8730
rect 7325 8678 7377 8730
rect 7389 8678 7441 8730
rect 7453 8678 7505 8730
rect 7517 8678 7569 8730
rect 7581 8678 7633 8730
rect 3976 8551 4028 8560
rect 3976 8517 3985 8551
rect 3985 8517 4019 8551
rect 4019 8517 4028 8551
rect 3976 8508 4028 8517
rect 4436 8440 4488 8492
rect 1766 8134 1818 8186
rect 1830 8134 1882 8186
rect 1894 8134 1946 8186
rect 1958 8134 2010 8186
rect 2022 8134 2074 8186
rect 3399 8134 3451 8186
rect 3463 8134 3515 8186
rect 3527 8134 3579 8186
rect 3591 8134 3643 8186
rect 3655 8134 3707 8186
rect 5032 8134 5084 8186
rect 5096 8134 5148 8186
rect 5160 8134 5212 8186
rect 5224 8134 5276 8186
rect 5288 8134 5340 8186
rect 6665 8134 6717 8186
rect 6729 8134 6781 8186
rect 6793 8134 6845 8186
rect 6857 8134 6909 8186
rect 6921 8134 6973 8186
rect 6184 7828 6236 7880
rect 7748 7828 7800 7880
rect 2426 7590 2478 7642
rect 2490 7590 2542 7642
rect 2554 7590 2606 7642
rect 2618 7590 2670 7642
rect 2682 7590 2734 7642
rect 4059 7590 4111 7642
rect 4123 7590 4175 7642
rect 4187 7590 4239 7642
rect 4251 7590 4303 7642
rect 4315 7590 4367 7642
rect 5692 7590 5744 7642
rect 5756 7590 5808 7642
rect 5820 7590 5872 7642
rect 5884 7590 5936 7642
rect 5948 7590 6000 7642
rect 7325 7590 7377 7642
rect 7389 7590 7441 7642
rect 7453 7590 7505 7642
rect 7517 7590 7569 7642
rect 7581 7590 7633 7642
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 3240 7420 3292 7472
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 3884 7352 3936 7404
rect 5540 7352 5592 7404
rect 6000 7352 6052 7404
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 6092 7259 6144 7268
rect 6092 7225 6101 7259
rect 6101 7225 6135 7259
rect 6135 7225 6144 7259
rect 6092 7216 6144 7225
rect 2228 7148 2280 7200
rect 3976 7148 4028 7200
rect 5724 7148 5776 7200
rect 6184 7148 6236 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 1766 7046 1818 7098
rect 1830 7046 1882 7098
rect 1894 7046 1946 7098
rect 1958 7046 2010 7098
rect 2022 7046 2074 7098
rect 3399 7046 3451 7098
rect 3463 7046 3515 7098
rect 3527 7046 3579 7098
rect 3591 7046 3643 7098
rect 3655 7046 3707 7098
rect 5032 7046 5084 7098
rect 5096 7046 5148 7098
rect 5160 7046 5212 7098
rect 5224 7046 5276 7098
rect 5288 7046 5340 7098
rect 6665 7046 6717 7098
rect 6729 7046 6781 7098
rect 6793 7046 6845 7098
rect 6857 7046 6909 7098
rect 6921 7046 6973 7098
rect 2136 6851 2188 6860
rect 2136 6817 2145 6851
rect 2145 6817 2179 6851
rect 2179 6817 2188 6851
rect 2136 6808 2188 6817
rect 3148 6808 3200 6860
rect 5816 6944 5868 6996
rect 5264 6876 5316 6928
rect 6644 6876 6696 6928
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2596 6740 2648 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 2136 6672 2188 6724
rect 2596 6647 2648 6656
rect 2596 6613 2605 6647
rect 2605 6613 2639 6647
rect 2639 6613 2648 6647
rect 2596 6604 2648 6613
rect 3332 6672 3384 6724
rect 3608 6672 3660 6724
rect 4620 6740 4672 6792
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 6092 6808 6144 6860
rect 6736 6740 6788 6792
rect 5448 6604 5500 6656
rect 6552 6715 6604 6724
rect 6552 6681 6561 6715
rect 6561 6681 6595 6715
rect 6595 6681 6604 6715
rect 6552 6672 6604 6681
rect 2426 6502 2478 6554
rect 2490 6502 2542 6554
rect 2554 6502 2606 6554
rect 2618 6502 2670 6554
rect 2682 6502 2734 6554
rect 4059 6502 4111 6554
rect 4123 6502 4175 6554
rect 4187 6502 4239 6554
rect 4251 6502 4303 6554
rect 4315 6502 4367 6554
rect 5692 6502 5744 6554
rect 5756 6502 5808 6554
rect 5820 6502 5872 6554
rect 5884 6502 5936 6554
rect 5948 6502 6000 6554
rect 7325 6502 7377 6554
rect 7389 6502 7441 6554
rect 7453 6502 7505 6554
rect 7517 6502 7569 6554
rect 7581 6502 7633 6554
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 5356 6400 5408 6452
rect 6552 6400 6604 6452
rect 6644 6400 6696 6452
rect 848 6264 900 6316
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 4528 6196 4580 6248
rect 3240 6128 3292 6180
rect 3884 6128 3936 6180
rect 5356 6264 5408 6316
rect 5724 6264 5776 6316
rect 6184 6264 6236 6316
rect 6000 6196 6052 6248
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 4804 6128 4856 6180
rect 5724 6128 5776 6180
rect 4620 6060 4672 6112
rect 6184 6060 6236 6112
rect 1766 5958 1818 6010
rect 1830 5958 1882 6010
rect 1894 5958 1946 6010
rect 1958 5958 2010 6010
rect 2022 5958 2074 6010
rect 3399 5958 3451 6010
rect 3463 5958 3515 6010
rect 3527 5958 3579 6010
rect 3591 5958 3643 6010
rect 3655 5958 3707 6010
rect 5032 5958 5084 6010
rect 5096 5958 5148 6010
rect 5160 5958 5212 6010
rect 5224 5958 5276 6010
rect 5288 5958 5340 6010
rect 6665 5958 6717 6010
rect 6729 5958 6781 6010
rect 6793 5958 6845 6010
rect 6857 5958 6909 6010
rect 6921 5958 6973 6010
rect 2136 5856 2188 5908
rect 5356 5788 5408 5840
rect 4436 5720 4488 5772
rect 4528 5652 4580 5704
rect 7748 5652 7800 5704
rect 2426 5414 2478 5466
rect 2490 5414 2542 5466
rect 2554 5414 2606 5466
rect 2618 5414 2670 5466
rect 2682 5414 2734 5466
rect 4059 5414 4111 5466
rect 4123 5414 4175 5466
rect 4187 5414 4239 5466
rect 4251 5414 4303 5466
rect 4315 5414 4367 5466
rect 5692 5414 5744 5466
rect 5756 5414 5808 5466
rect 5820 5414 5872 5466
rect 5884 5414 5936 5466
rect 5948 5414 6000 5466
rect 7325 5414 7377 5466
rect 7389 5414 7441 5466
rect 7453 5414 7505 5466
rect 7517 5414 7569 5466
rect 7581 5414 7633 5466
rect 4436 5312 4488 5364
rect 4804 5355 4856 5364
rect 4804 5321 4813 5355
rect 4813 5321 4847 5355
rect 4847 5321 4856 5355
rect 4804 5312 4856 5321
rect 6092 5312 6144 5364
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 4804 5108 4856 5160
rect 6092 5176 6144 5228
rect 6276 5176 6328 5228
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 4160 5040 4212 5092
rect 6184 5083 6236 5092
rect 6184 5049 6193 5083
rect 6193 5049 6227 5083
rect 6227 5049 6236 5083
rect 6184 5040 6236 5049
rect 6276 4972 6328 5024
rect 1766 4870 1818 4922
rect 1830 4870 1882 4922
rect 1894 4870 1946 4922
rect 1958 4870 2010 4922
rect 2022 4870 2074 4922
rect 3399 4870 3451 4922
rect 3463 4870 3515 4922
rect 3527 4870 3579 4922
rect 3591 4870 3643 4922
rect 3655 4870 3707 4922
rect 5032 4870 5084 4922
rect 5096 4870 5148 4922
rect 5160 4870 5212 4922
rect 5224 4870 5276 4922
rect 5288 4870 5340 4922
rect 6665 4870 6717 4922
rect 6729 4870 6781 4922
rect 6793 4870 6845 4922
rect 6857 4870 6909 4922
rect 6921 4870 6973 4922
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 4896 4768 4948 4820
rect 5356 4768 5408 4820
rect 4160 4743 4212 4752
rect 4160 4709 4169 4743
rect 4169 4709 4203 4743
rect 4203 4709 4212 4743
rect 4160 4700 4212 4709
rect 4528 4700 4580 4752
rect 5448 4564 5500 4616
rect 7748 4564 7800 4616
rect 6092 4496 6144 4548
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 2426 4326 2478 4378
rect 2490 4326 2542 4378
rect 2554 4326 2606 4378
rect 2618 4326 2670 4378
rect 2682 4326 2734 4378
rect 4059 4326 4111 4378
rect 4123 4326 4175 4378
rect 4187 4326 4239 4378
rect 4251 4326 4303 4378
rect 4315 4326 4367 4378
rect 5692 4326 5744 4378
rect 5756 4326 5808 4378
rect 5820 4326 5872 4378
rect 5884 4326 5936 4378
rect 5948 4326 6000 4378
rect 7325 4326 7377 4378
rect 7389 4326 7441 4378
rect 7453 4326 7505 4378
rect 7517 4326 7569 4378
rect 7581 4326 7633 4378
rect 2780 4088 2832 4140
rect 2964 4088 3016 4140
rect 6092 4156 6144 4208
rect 6184 4088 6236 4140
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 1766 3782 1818 3834
rect 1830 3782 1882 3834
rect 1894 3782 1946 3834
rect 1958 3782 2010 3834
rect 2022 3782 2074 3834
rect 3399 3782 3451 3834
rect 3463 3782 3515 3834
rect 3527 3782 3579 3834
rect 3591 3782 3643 3834
rect 3655 3782 3707 3834
rect 5032 3782 5084 3834
rect 5096 3782 5148 3834
rect 5160 3782 5212 3834
rect 5224 3782 5276 3834
rect 5288 3782 5340 3834
rect 6665 3782 6717 3834
rect 6729 3782 6781 3834
rect 6793 3782 6845 3834
rect 6857 3782 6909 3834
rect 6921 3782 6973 3834
rect 2964 3680 3016 3732
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 3148 3544 3200 3596
rect 3884 3544 3936 3596
rect 5540 3680 5592 3732
rect 6184 3723 6236 3732
rect 6184 3689 6193 3723
rect 6193 3689 6227 3723
rect 6227 3689 6236 3723
rect 6184 3680 6236 3689
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 2872 3476 2924 3528
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 4620 3476 4672 3528
rect 6092 3476 6144 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 2872 3340 2924 3392
rect 4436 3408 4488 3460
rect 5356 3408 5408 3460
rect 4528 3383 4580 3392
rect 4528 3349 4537 3383
rect 4537 3349 4571 3383
rect 4571 3349 4580 3383
rect 4528 3340 4580 3349
rect 5448 3340 5500 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 2426 3238 2478 3290
rect 2490 3238 2542 3290
rect 2554 3238 2606 3290
rect 2618 3238 2670 3290
rect 2682 3238 2734 3290
rect 4059 3238 4111 3290
rect 4123 3238 4175 3290
rect 4187 3238 4239 3290
rect 4251 3238 4303 3290
rect 4315 3238 4367 3290
rect 5692 3238 5744 3290
rect 5756 3238 5808 3290
rect 5820 3238 5872 3290
rect 5884 3238 5936 3290
rect 5948 3238 6000 3290
rect 7325 3238 7377 3290
rect 7389 3238 7441 3290
rect 7453 3238 7505 3290
rect 7517 3238 7569 3290
rect 7581 3238 7633 3290
rect 2780 3136 2832 3188
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3792 3136 3844 3188
rect 7012 3136 7064 3188
rect 2320 3068 2372 3120
rect 2872 3068 2924 3120
rect 2136 3000 2188 3052
rect 2688 3000 2740 3052
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 4436 3000 4488 3052
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6092 3000 6144 3052
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 6184 2864 6236 2916
rect 1766 2694 1818 2746
rect 1830 2694 1882 2746
rect 1894 2694 1946 2746
rect 1958 2694 2010 2746
rect 2022 2694 2074 2746
rect 3399 2694 3451 2746
rect 3463 2694 3515 2746
rect 3527 2694 3579 2746
rect 3591 2694 3643 2746
rect 3655 2694 3707 2746
rect 5032 2694 5084 2746
rect 5096 2694 5148 2746
rect 5160 2694 5212 2746
rect 5224 2694 5276 2746
rect 5288 2694 5340 2746
rect 6665 2694 6717 2746
rect 6729 2694 6781 2746
rect 6793 2694 6845 2746
rect 6857 2694 6909 2746
rect 6921 2694 6973 2746
rect 2688 2635 2740 2644
rect 2688 2601 2697 2635
rect 2697 2601 2731 2635
rect 2731 2601 2740 2635
rect 2688 2592 2740 2601
rect 2780 2592 2832 2644
rect 2320 2388 2372 2440
rect 3240 2388 3292 2440
rect 4528 2388 4580 2440
rect 3884 2252 3936 2304
rect 2426 2150 2478 2202
rect 2490 2150 2542 2202
rect 2554 2150 2606 2202
rect 2618 2150 2670 2202
rect 2682 2150 2734 2202
rect 4059 2150 4111 2202
rect 4123 2150 4175 2202
rect 4187 2150 4239 2202
rect 4251 2150 4303 2202
rect 4315 2150 4367 2202
rect 5692 2150 5744 2202
rect 5756 2150 5808 2202
rect 5820 2150 5872 2202
rect 5884 2150 5936 2202
rect 5948 2150 6000 2202
rect 7325 2150 7377 2202
rect 7389 2150 7441 2202
rect 7453 2150 7505 2202
rect 7517 2150 7569 2202
rect 7581 2150 7633 2202
<< metal2 >>
rect 3882 10282 3938 10963
rect 3882 10254 4016 10282
rect 3882 10163 3938 10254
rect 2426 8732 2734 8741
rect 2426 8730 2432 8732
rect 2488 8730 2512 8732
rect 2568 8730 2592 8732
rect 2648 8730 2672 8732
rect 2728 8730 2734 8732
rect 2488 8678 2490 8730
rect 2670 8678 2672 8730
rect 2426 8676 2432 8678
rect 2488 8676 2512 8678
rect 2568 8676 2592 8678
rect 2648 8676 2672 8678
rect 2728 8676 2734 8678
rect 2426 8667 2734 8676
rect 3988 8566 4016 10254
rect 4059 8732 4367 8741
rect 4059 8730 4065 8732
rect 4121 8730 4145 8732
rect 4201 8730 4225 8732
rect 4281 8730 4305 8732
rect 4361 8730 4367 8732
rect 4121 8678 4123 8730
rect 4303 8678 4305 8730
rect 4059 8676 4065 8678
rect 4121 8676 4145 8678
rect 4201 8676 4225 8678
rect 4281 8676 4305 8678
rect 4361 8676 4367 8678
rect 4059 8667 4367 8676
rect 5692 8732 6000 8741
rect 5692 8730 5698 8732
rect 5754 8730 5778 8732
rect 5834 8730 5858 8732
rect 5914 8730 5938 8732
rect 5994 8730 6000 8732
rect 5754 8678 5756 8730
rect 5936 8678 5938 8730
rect 5692 8676 5698 8678
rect 5754 8676 5778 8678
rect 5834 8676 5858 8678
rect 5914 8676 5938 8678
rect 5994 8676 6000 8678
rect 5692 8667 6000 8676
rect 7325 8732 7633 8741
rect 7325 8730 7331 8732
rect 7387 8730 7411 8732
rect 7467 8730 7491 8732
rect 7547 8730 7571 8732
rect 7627 8730 7633 8732
rect 7387 8678 7389 8730
rect 7569 8678 7571 8730
rect 7325 8676 7331 8678
rect 7387 8676 7411 8678
rect 7467 8676 7491 8678
rect 7547 8676 7571 8678
rect 7627 8676 7633 8678
rect 7325 8667 7633 8676
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 1766 8188 2074 8197
rect 1766 8186 1772 8188
rect 1828 8186 1852 8188
rect 1908 8186 1932 8188
rect 1988 8186 2012 8188
rect 2068 8186 2074 8188
rect 1828 8134 1830 8186
rect 2010 8134 2012 8186
rect 1766 8132 1772 8134
rect 1828 8132 1852 8134
rect 1908 8132 1932 8134
rect 1988 8132 2012 8134
rect 2068 8132 2074 8134
rect 1766 8123 2074 8132
rect 3399 8188 3707 8197
rect 3399 8186 3405 8188
rect 3461 8186 3485 8188
rect 3541 8186 3565 8188
rect 3621 8186 3645 8188
rect 3701 8186 3707 8188
rect 3461 8134 3463 8186
rect 3643 8134 3645 8186
rect 3399 8132 3405 8134
rect 3461 8132 3485 8134
rect 3541 8132 3565 8134
rect 3621 8132 3645 8134
rect 3701 8132 3707 8134
rect 3399 8123 3707 8132
rect 2426 7644 2734 7653
rect 2426 7642 2432 7644
rect 2488 7642 2512 7644
rect 2568 7642 2592 7644
rect 2648 7642 2672 7644
rect 2728 7642 2734 7644
rect 2488 7590 2490 7642
rect 2670 7590 2672 7642
rect 2426 7588 2432 7590
rect 2488 7588 2512 7590
rect 2568 7588 2592 7590
rect 2648 7588 2672 7590
rect 2728 7588 2734 7590
rect 2426 7579 2734 7588
rect 4059 7644 4367 7653
rect 4059 7642 4065 7644
rect 4121 7642 4145 7644
rect 4201 7642 4225 7644
rect 4281 7642 4305 7644
rect 4361 7642 4367 7644
rect 4121 7590 4123 7642
rect 4303 7590 4305 7642
rect 4059 7588 4065 7590
rect 4121 7588 4145 7590
rect 4201 7588 4225 7590
rect 4281 7588 4305 7590
rect 4361 7588 4367 7590
rect 4059 7579 4367 7588
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 1766 7100 2074 7109
rect 1766 7098 1772 7100
rect 1828 7098 1852 7100
rect 1908 7098 1932 7100
rect 1988 7098 2012 7100
rect 2068 7098 2074 7100
rect 1828 7046 1830 7098
rect 2010 7046 2012 7098
rect 1766 7044 1772 7046
rect 1828 7044 1852 7046
rect 1908 7044 1932 7046
rect 1988 7044 2012 7046
rect 2068 7044 2074 7046
rect 1766 7035 2074 7044
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2148 6730 2176 6802
rect 2240 6798 2268 7142
rect 2608 6798 2636 7278
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1766 6012 2074 6021
rect 1766 6010 1772 6012
rect 1828 6010 1852 6012
rect 1908 6010 1932 6012
rect 1988 6010 2012 6012
rect 2068 6010 2074 6012
rect 1828 5958 1830 6010
rect 2010 5958 2012 6010
rect 1766 5956 1772 5958
rect 1828 5956 1852 5958
rect 1908 5956 1932 5958
rect 1988 5956 2012 5958
rect 2068 5956 2074 5958
rect 1766 5947 2074 5956
rect 2148 5914 2176 6666
rect 2608 6662 2636 6734
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2426 6556 2734 6565
rect 2426 6554 2432 6556
rect 2488 6554 2512 6556
rect 2568 6554 2592 6556
rect 2648 6554 2672 6556
rect 2728 6554 2734 6556
rect 2488 6502 2490 6554
rect 2670 6502 2672 6554
rect 2426 6500 2432 6502
rect 2488 6500 2512 6502
rect 2568 6500 2592 6502
rect 2648 6500 2672 6502
rect 2728 6500 2734 6502
rect 2426 6491 2734 6500
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2426 5468 2734 5477
rect 2426 5466 2432 5468
rect 2488 5466 2512 5468
rect 2568 5466 2592 5468
rect 2648 5466 2672 5468
rect 2728 5466 2734 5468
rect 2488 5414 2490 5466
rect 2670 5414 2672 5466
rect 2426 5412 2432 5414
rect 2488 5412 2512 5414
rect 2568 5412 2592 5414
rect 2648 5412 2672 5414
rect 2728 5412 2734 5414
rect 2426 5403 2734 5412
rect 1766 4924 2074 4933
rect 1766 4922 1772 4924
rect 1828 4922 1852 4924
rect 1908 4922 1932 4924
rect 1988 4922 2012 4924
rect 2068 4922 2074 4924
rect 1828 4870 1830 4922
rect 2010 4870 2012 4922
rect 1766 4868 1772 4870
rect 1828 4868 1852 4870
rect 1908 4868 1932 4870
rect 1988 4868 2012 4870
rect 2068 4868 2074 4870
rect 1766 4859 2074 4868
rect 2426 4380 2734 4389
rect 2426 4378 2432 4380
rect 2488 4378 2512 4380
rect 2568 4378 2592 4380
rect 2648 4378 2672 4380
rect 2728 4378 2734 4380
rect 2488 4326 2490 4378
rect 2670 4326 2672 4378
rect 2426 4324 2432 4326
rect 2488 4324 2512 4326
rect 2568 4324 2592 4326
rect 2648 4324 2672 4326
rect 2728 4324 2734 4326
rect 2426 4315 2734 4324
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 1766 3836 2074 3845
rect 1766 3834 1772 3836
rect 1828 3834 1852 3836
rect 1908 3834 1932 3836
rect 1988 3834 2012 3836
rect 2068 3834 2074 3836
rect 1828 3782 1830 3834
rect 2010 3782 2012 3834
rect 1766 3780 1772 3782
rect 1828 3780 1852 3782
rect 1908 3780 1932 3782
rect 1988 3780 2012 3782
rect 2068 3780 2074 3782
rect 1766 3771 2074 3780
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2148 3058 2176 3470
rect 2332 3126 2360 3470
rect 2792 3346 2820 4082
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3534 2912 3878
rect 2976 3738 3004 4082
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2872 3392 2924 3398
rect 2792 3340 2872 3346
rect 2792 3334 2924 3340
rect 2792 3318 2912 3334
rect 2426 3292 2734 3301
rect 2426 3290 2432 3292
rect 2488 3290 2512 3292
rect 2568 3290 2592 3292
rect 2648 3290 2672 3292
rect 2728 3290 2734 3292
rect 2488 3238 2490 3290
rect 2670 3238 2672 3290
rect 2426 3236 2432 3238
rect 2488 3236 2512 3238
rect 2568 3236 2592 3238
rect 2648 3236 2672 3238
rect 2728 3236 2734 3238
rect 2426 3227 2734 3236
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2792 3058 2820 3130
rect 2884 3126 2912 3318
rect 2976 3194 3004 3674
rect 3160 3602 3188 6802
rect 3252 6746 3280 7414
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3399 7100 3707 7109
rect 3399 7098 3405 7100
rect 3461 7098 3485 7100
rect 3541 7098 3565 7100
rect 3621 7098 3645 7100
rect 3701 7098 3707 7100
rect 3461 7046 3463 7098
rect 3643 7046 3645 7098
rect 3399 7044 3405 7046
rect 3461 7044 3485 7046
rect 3541 7044 3565 7046
rect 3621 7044 3645 7046
rect 3701 7044 3707 7046
rect 3399 7035 3707 7044
rect 3792 6792 3844 6798
rect 3252 6730 3372 6746
rect 3792 6734 3844 6740
rect 3252 6724 3384 6730
rect 3252 6718 3332 6724
rect 3332 6666 3384 6672
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3620 6322 3648 6666
rect 3804 6458 3832 6734
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3252 6186 3280 6258
rect 3896 6186 3924 7346
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6798 4016 7142
rect 4448 6866 4476 8434
rect 5032 8188 5340 8197
rect 5032 8186 5038 8188
rect 5094 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5340 8188
rect 5094 8134 5096 8186
rect 5276 8134 5278 8186
rect 5032 8132 5038 8134
rect 5094 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5340 8134
rect 5032 8123 5340 8132
rect 6665 8188 6973 8197
rect 6665 8186 6671 8188
rect 6727 8186 6751 8188
rect 6807 8186 6831 8188
rect 6887 8186 6911 8188
rect 6967 8186 6973 8188
rect 6727 8134 6729 8186
rect 6909 8134 6911 8186
rect 6665 8132 6671 8134
rect 6727 8132 6751 8134
rect 6807 8132 6831 8134
rect 6887 8132 6911 8134
rect 6967 8132 6973 8134
rect 6665 8123 6973 8132
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 5692 7644 6000 7653
rect 5692 7642 5698 7644
rect 5754 7642 5778 7644
rect 5834 7642 5858 7644
rect 5914 7642 5938 7644
rect 5994 7642 6000 7644
rect 5754 7590 5756 7642
rect 5936 7590 5938 7642
rect 5692 7588 5698 7590
rect 5754 7588 5778 7590
rect 5834 7588 5858 7590
rect 5914 7588 5938 7590
rect 5994 7588 6000 7590
rect 5692 7579 6000 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5032 7100 5340 7109
rect 5032 7098 5038 7100
rect 5094 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5340 7100
rect 5094 7046 5096 7098
rect 5276 7046 5278 7098
rect 5032 7044 5038 7046
rect 5094 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5340 7046
rect 5032 7035 5340 7044
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 5276 6798 5304 6870
rect 3976 6792 4028 6798
rect 4620 6792 4672 6798
rect 3976 6734 4028 6740
rect 4618 6760 4620 6769
rect 5264 6792 5316 6798
rect 4672 6760 4674 6769
rect 5264 6734 5316 6740
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 4618 6695 4674 6704
rect 4059 6556 4367 6565
rect 4059 6554 4065 6556
rect 4121 6554 4145 6556
rect 4201 6554 4225 6556
rect 4281 6554 4305 6556
rect 4361 6554 4367 6556
rect 4121 6502 4123 6554
rect 4303 6502 4305 6554
rect 4059 6500 4065 6502
rect 4121 6500 4145 6502
rect 4201 6500 4225 6502
rect 4281 6500 4305 6502
rect 4361 6500 4367 6502
rect 4059 6491 4367 6500
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3399 6012 3707 6021
rect 3399 6010 3405 6012
rect 3461 6010 3485 6012
rect 3541 6010 3565 6012
rect 3621 6010 3645 6012
rect 3701 6010 3707 6012
rect 3461 5958 3463 6010
rect 3643 5958 3645 6010
rect 3399 5956 3405 5958
rect 3461 5956 3485 5958
rect 3541 5956 3565 5958
rect 3621 5956 3645 5958
rect 3701 5956 3707 5958
rect 3399 5947 3707 5956
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4059 5468 4367 5477
rect 4059 5466 4065 5468
rect 4121 5466 4145 5468
rect 4201 5466 4225 5468
rect 4281 5466 4305 5468
rect 4361 5466 4367 5468
rect 4121 5414 4123 5466
rect 4303 5414 4305 5466
rect 4059 5412 4065 5414
rect 4121 5412 4145 5414
rect 4201 5412 4225 5414
rect 4281 5412 4305 5414
rect 4361 5412 4367 5414
rect 4059 5403 4367 5412
rect 4448 5370 4476 5714
rect 4540 5710 4568 6190
rect 4632 6118 4660 6695
rect 5368 6458 5396 6734
rect 5448 6656 5500 6662
rect 5552 6644 5580 7346
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 6798 5764 7142
rect 5828 7002 5856 7278
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 6012 6866 6040 7346
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6104 6866 6132 7210
rect 6196 7206 6224 7822
rect 7325 7644 7633 7653
rect 7325 7642 7331 7644
rect 7387 7642 7411 7644
rect 7467 7642 7491 7644
rect 7547 7642 7571 7644
rect 7627 7642 7633 7644
rect 7387 7590 7389 7642
rect 7569 7590 7571 7642
rect 7325 7588 7331 7590
rect 7387 7588 7411 7590
rect 7467 7588 7491 7590
rect 7547 7588 7571 7590
rect 7627 7588 7633 7590
rect 7325 7579 7633 7588
rect 7760 7585 7788 7822
rect 7746 7576 7802 7585
rect 7746 7511 7802 7520
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5632 6792 5684 6798
rect 5630 6760 5632 6769
rect 5724 6792 5776 6798
rect 5684 6760 5686 6769
rect 5724 6734 5776 6740
rect 5630 6695 5686 6704
rect 5500 6616 5580 6644
rect 5448 6598 5500 6604
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3399 4924 3707 4933
rect 3399 4922 3405 4924
rect 3461 4922 3485 4924
rect 3541 4922 3565 4924
rect 3621 4922 3645 4924
rect 3701 4922 3707 4924
rect 3461 4870 3463 4922
rect 3643 4870 3645 4922
rect 3399 4868 3405 4870
rect 3461 4868 3485 4870
rect 3541 4868 3565 4870
rect 3621 4868 3645 4870
rect 3701 4868 3707 4870
rect 3399 4859 3707 4868
rect 4172 4758 4200 5034
rect 4540 4758 4568 5646
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3399 3836 3707 3845
rect 3399 3834 3405 3836
rect 3461 3834 3485 3836
rect 3541 3834 3565 3836
rect 3621 3834 3645 3836
rect 3701 3834 3707 3836
rect 3461 3782 3463 3834
rect 3643 3782 3645 3834
rect 3399 3780 3405 3782
rect 3461 3780 3485 3782
rect 3541 3780 3565 3782
rect 3621 3780 3645 3782
rect 3701 3780 3707 3782
rect 3399 3771 3707 3780
rect 3896 3602 3924 4422
rect 4059 4380 4367 4389
rect 4059 4378 4065 4380
rect 4121 4378 4145 4380
rect 4201 4378 4225 4380
rect 4281 4378 4305 4380
rect 4361 4378 4367 4380
rect 4121 4326 4123 4378
rect 4303 4326 4305 4378
rect 4059 4324 4065 4326
rect 4121 4324 4145 4326
rect 4201 4324 4225 4326
rect 4281 4324 4305 4326
rect 4361 4324 4367 4326
rect 4059 4315 4367 4324
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 4632 3534 4660 6054
rect 4816 5370 4844 6122
rect 5032 6012 5340 6021
rect 5032 6010 5038 6012
rect 5094 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5340 6012
rect 5094 5958 5096 6010
rect 5276 5958 5278 6010
rect 5032 5956 5038 5958
rect 5094 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5340 5958
rect 5032 5947 5340 5956
rect 5368 5846 5396 6258
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4816 4826 4844 5102
rect 4908 4826 4936 5170
rect 5368 4978 5396 5782
rect 5368 4950 5488 4978
rect 5032 4924 5340 4933
rect 5032 4922 5038 4924
rect 5094 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5340 4924
rect 5094 4870 5096 4922
rect 5276 4870 5278 4922
rect 5032 4868 5038 4870
rect 5094 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5340 4870
rect 5032 4859 5340 4868
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5032 3836 5340 3845
rect 5032 3834 5038 3836
rect 5094 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5340 3836
rect 5094 3782 5096 3834
rect 5276 3782 5278 3834
rect 5032 3780 5038 3782
rect 5094 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5340 3782
rect 5032 3771 5340 3780
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 3804 3194 3832 3470
rect 5368 3466 5396 4762
rect 5460 4622 5488 4950
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5552 3738 5580 6616
rect 5692 6556 6000 6565
rect 5692 6554 5698 6556
rect 5754 6554 5778 6556
rect 5834 6554 5858 6556
rect 5914 6554 5938 6556
rect 5994 6554 6000 6556
rect 5754 6502 5756 6554
rect 5936 6502 5938 6554
rect 5692 6500 5698 6502
rect 5754 6500 5778 6502
rect 5834 6500 5858 6502
rect 5914 6500 5938 6502
rect 5994 6500 6000 6502
rect 5692 6491 6000 6500
rect 6196 6474 6224 7142
rect 6665 7100 6973 7109
rect 6665 7098 6671 7100
rect 6727 7098 6751 7100
rect 6807 7098 6831 7100
rect 6887 7098 6911 7100
rect 6967 7098 6973 7100
rect 6727 7046 6729 7098
rect 6909 7046 6911 7098
rect 6665 7044 6671 7046
rect 6727 7044 6751 7046
rect 6807 7044 6831 7046
rect 6887 7044 6911 7046
rect 6967 7044 6973 7046
rect 6665 7035 6973 7044
rect 6644 6928 6696 6934
rect 7208 6905 7236 7142
rect 6644 6870 6696 6876
rect 7194 6896 7250 6905
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6104 6446 6316 6474
rect 6564 6458 6592 6666
rect 6656 6458 6684 6870
rect 7194 6831 7250 6840
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 5722 6352 5778 6361
rect 6104 6338 6132 6446
rect 5722 6287 5724 6296
rect 5776 6287 5778 6296
rect 6012 6310 6132 6338
rect 6184 6316 6236 6322
rect 5724 6258 5776 6264
rect 5736 6186 5764 6258
rect 6012 6254 6040 6310
rect 6184 6258 6236 6264
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5692 5468 6000 5477
rect 5692 5466 5698 5468
rect 5754 5466 5778 5468
rect 5834 5466 5858 5468
rect 5914 5466 5938 5468
rect 5994 5466 6000 5468
rect 5754 5414 5756 5466
rect 5936 5414 5938 5466
rect 5692 5412 5698 5414
rect 5754 5412 5778 5414
rect 5834 5412 5858 5414
rect 5914 5412 5938 5414
rect 5994 5412 6000 5414
rect 5692 5403 6000 5412
rect 6104 5370 6132 6190
rect 6196 6118 6224 6258
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6104 4554 6132 5170
rect 6196 5098 6224 6054
rect 6288 5234 6316 6446
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6748 6361 6776 6734
rect 7325 6556 7633 6565
rect 7325 6554 7331 6556
rect 7387 6554 7411 6556
rect 7467 6554 7491 6556
rect 7547 6554 7571 6556
rect 7627 6554 7633 6556
rect 7387 6502 7389 6554
rect 7569 6502 7571 6554
rect 7325 6500 7331 6502
rect 7387 6500 7411 6502
rect 7467 6500 7491 6502
rect 7547 6500 7571 6502
rect 7627 6500 7633 6502
rect 7325 6491 7633 6500
rect 6734 6352 6790 6361
rect 6734 6287 6790 6296
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7300 6225 7328 6258
rect 7286 6216 7342 6225
rect 7286 6151 7342 6160
rect 6665 6012 6973 6021
rect 6665 6010 6671 6012
rect 6727 6010 6751 6012
rect 6807 6010 6831 6012
rect 6887 6010 6911 6012
rect 6967 6010 6973 6012
rect 6727 5958 6729 6010
rect 6909 5958 6911 6010
rect 6665 5956 6671 5958
rect 6727 5956 6751 5958
rect 6807 5956 6831 5958
rect 6887 5956 6911 5958
rect 6967 5956 6973 5958
rect 6665 5947 6973 5956
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7760 5545 7788 5646
rect 7746 5536 7802 5545
rect 7325 5468 7633 5477
rect 7746 5471 7802 5480
rect 7325 5466 7331 5468
rect 7387 5466 7411 5468
rect 7467 5466 7491 5468
rect 7547 5466 7571 5468
rect 7627 5466 7633 5468
rect 7387 5414 7389 5466
rect 7569 5414 7571 5466
rect 7325 5412 7331 5414
rect 7387 5412 7411 5414
rect 7467 5412 7491 5414
rect 7547 5412 7571 5414
rect 7627 5412 7633 5414
rect 7325 5403 7633 5412
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6288 5030 6316 5170
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6665 4924 6973 4933
rect 6665 4922 6671 4924
rect 6727 4922 6751 4924
rect 6807 4922 6831 4924
rect 6887 4922 6911 4924
rect 6967 4922 6973 4924
rect 6727 4870 6729 4922
rect 6909 4870 6911 4922
rect 6665 4868 6671 4870
rect 6727 4868 6751 4870
rect 6807 4868 6831 4870
rect 6887 4868 6911 4870
rect 6967 4868 6973 4870
rect 6665 4859 6973 4868
rect 7208 4865 7236 5170
rect 7194 4856 7250 4865
rect 7194 4791 7250 4800
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 5692 4380 6000 4389
rect 5692 4378 5698 4380
rect 5754 4378 5778 4380
rect 5834 4378 5858 4380
rect 5914 4378 5938 4380
rect 5994 4378 6000 4380
rect 5754 4326 5756 4378
rect 5936 4326 5938 4378
rect 5692 4324 5698 4326
rect 5754 4324 5778 4326
rect 5834 4324 5858 4326
rect 5914 4324 5938 4326
rect 5994 4324 6000 4326
rect 5692 4315 6000 4324
rect 6104 4214 6132 4490
rect 7325 4380 7633 4389
rect 7325 4378 7331 4380
rect 7387 4378 7411 4380
rect 7467 4378 7491 4380
rect 7547 4378 7571 4380
rect 7627 4378 7633 4380
rect 7387 4326 7389 4378
rect 7569 4326 7571 4378
rect 7325 4324 7331 4326
rect 7387 4324 7411 4326
rect 7467 4324 7491 4326
rect 7547 4324 7571 4326
rect 7627 4324 7633 4326
rect 7325 4315 7633 4324
rect 6092 4208 6144 4214
rect 7760 4185 7788 4558
rect 6092 4150 6144 4156
rect 7746 4176 7802 4185
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5736 3602 5764 3878
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 6104 3534 6132 4150
rect 6184 4140 6236 4146
rect 7746 4111 7802 4120
rect 6184 4082 6236 4088
rect 6196 3738 6224 4082
rect 6665 3836 6973 3845
rect 6665 3834 6671 3836
rect 6727 3834 6751 3836
rect 6807 3834 6831 3836
rect 6887 3834 6911 3836
rect 6967 3834 6973 3836
rect 6727 3782 6729 3834
rect 6909 3782 6911 3834
rect 6665 3780 6671 3782
rect 6727 3780 6751 3782
rect 6807 3780 6831 3782
rect 6887 3780 6911 3782
rect 6967 3780 6973 3782
rect 6665 3771 6973 3780
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 4059 3292 4367 3301
rect 4059 3290 4065 3292
rect 4121 3290 4145 3292
rect 4201 3290 4225 3292
rect 4281 3290 4305 3292
rect 4361 3290 4367 3292
rect 4121 3238 4123 3290
rect 4303 3238 4305 3290
rect 4059 3236 4065 3238
rect 4121 3236 4145 3238
rect 4201 3236 4225 3238
rect 4281 3236 4305 3238
rect 4361 3236 4367 3238
rect 4059 3227 4367 3236
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 4448 3058 4476 3402
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 1766 2748 2074 2757
rect 1766 2746 1772 2748
rect 1828 2746 1852 2748
rect 1908 2746 1932 2748
rect 1988 2746 2012 2748
rect 2068 2746 2074 2748
rect 1828 2694 1830 2746
rect 2010 2694 2012 2746
rect 1766 2692 1772 2694
rect 1828 2692 1852 2694
rect 1908 2692 1932 2694
rect 1988 2692 2012 2694
rect 2068 2692 2074 2694
rect 1766 2683 2074 2692
rect 2700 2650 2728 2994
rect 2792 2650 2820 2994
rect 3399 2748 3707 2757
rect 3399 2746 3405 2748
rect 3461 2746 3485 2748
rect 3541 2746 3565 2748
rect 3621 2746 3645 2748
rect 3701 2746 3707 2748
rect 3461 2694 3463 2746
rect 3643 2694 3645 2746
rect 3399 2692 3405 2694
rect 3461 2692 3485 2694
rect 3541 2692 3565 2694
rect 3621 2692 3645 2694
rect 3701 2692 3707 2694
rect 3399 2683 3707 2692
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 4540 2446 4568 3334
rect 5460 3058 5488 3334
rect 5692 3292 6000 3301
rect 5692 3290 5698 3292
rect 5754 3290 5778 3292
rect 5834 3290 5858 3292
rect 5914 3290 5938 3292
rect 5994 3290 6000 3292
rect 5754 3238 5756 3290
rect 5936 3238 5938 3290
rect 5692 3236 5698 3238
rect 5754 3236 5778 3238
rect 5834 3236 5858 3238
rect 5914 3236 5938 3238
rect 5994 3236 6000 3238
rect 5692 3227 6000 3236
rect 6104 3058 6132 3470
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6196 2922 6224 3674
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7194 3496 7250 3505
rect 7024 3194 7052 3470
rect 7194 3431 7250 3440
rect 7208 3398 7236 3431
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7325 3292 7633 3301
rect 7325 3290 7331 3292
rect 7387 3290 7411 3292
rect 7467 3290 7491 3292
rect 7547 3290 7571 3292
rect 7627 3290 7633 3292
rect 7387 3238 7389 3290
rect 7569 3238 7571 3290
rect 7325 3236 7331 3238
rect 7387 3236 7411 3238
rect 7467 3236 7491 3238
rect 7547 3236 7571 3238
rect 7627 3236 7633 3238
rect 7325 3227 7633 3236
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 7300 2825 7328 2994
rect 7286 2816 7342 2825
rect 5032 2748 5340 2757
rect 5032 2746 5038 2748
rect 5094 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5340 2748
rect 5094 2694 5096 2746
rect 5276 2694 5278 2746
rect 5032 2692 5038 2694
rect 5094 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5340 2694
rect 5032 2683 5340 2692
rect 6665 2748 6973 2757
rect 7286 2751 7342 2760
rect 6665 2746 6671 2748
rect 6727 2746 6751 2748
rect 6807 2746 6831 2748
rect 6887 2746 6911 2748
rect 6967 2746 6973 2748
rect 6727 2694 6729 2746
rect 6909 2694 6911 2746
rect 6665 2692 6671 2694
rect 6727 2692 6751 2694
rect 6807 2692 6831 2694
rect 6887 2692 6911 2694
rect 6967 2692 6973 2694
rect 6665 2683 6973 2692
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 2332 762 2360 2382
rect 2426 2204 2734 2213
rect 2426 2202 2432 2204
rect 2488 2202 2512 2204
rect 2568 2202 2592 2204
rect 2648 2202 2672 2204
rect 2728 2202 2734 2204
rect 2488 2150 2490 2202
rect 2670 2150 2672 2202
rect 2426 2148 2432 2150
rect 2488 2148 2512 2150
rect 2568 2148 2592 2150
rect 2648 2148 2672 2150
rect 2728 2148 2734 2150
rect 2426 2139 2734 2148
rect 2516 870 2636 898
rect 2516 762 2544 870
rect 2608 800 2636 870
rect 3252 800 3280 2382
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 800 3924 2246
rect 4059 2204 4367 2213
rect 4059 2202 4065 2204
rect 4121 2202 4145 2204
rect 4201 2202 4225 2204
rect 4281 2202 4305 2204
rect 4361 2202 4367 2204
rect 4121 2150 4123 2202
rect 4303 2150 4305 2202
rect 4059 2148 4065 2150
rect 4121 2148 4145 2150
rect 4201 2148 4225 2150
rect 4281 2148 4305 2150
rect 4361 2148 4367 2150
rect 4059 2139 4367 2148
rect 5692 2204 6000 2213
rect 5692 2202 5698 2204
rect 5754 2202 5778 2204
rect 5834 2202 5858 2204
rect 5914 2202 5938 2204
rect 5994 2202 6000 2204
rect 5754 2150 5756 2202
rect 5936 2150 5938 2202
rect 5692 2148 5698 2150
rect 5754 2148 5778 2150
rect 5834 2148 5858 2150
rect 5914 2148 5938 2150
rect 5994 2148 6000 2150
rect 5692 2139 6000 2148
rect 7325 2204 7633 2213
rect 7325 2202 7331 2204
rect 7387 2202 7411 2204
rect 7467 2202 7491 2204
rect 7547 2202 7571 2204
rect 7627 2202 7633 2204
rect 7387 2150 7389 2202
rect 7569 2150 7571 2202
rect 7325 2148 7331 2150
rect 7387 2148 7411 2150
rect 7467 2148 7491 2150
rect 7547 2148 7571 2150
rect 7627 2148 7633 2150
rect 7325 2139 7633 2148
rect 2332 734 2544 762
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
<< via2 >>
rect 2432 8730 2488 8732
rect 2512 8730 2568 8732
rect 2592 8730 2648 8732
rect 2672 8730 2728 8732
rect 2432 8678 2478 8730
rect 2478 8678 2488 8730
rect 2512 8678 2542 8730
rect 2542 8678 2554 8730
rect 2554 8678 2568 8730
rect 2592 8678 2606 8730
rect 2606 8678 2618 8730
rect 2618 8678 2648 8730
rect 2672 8678 2682 8730
rect 2682 8678 2728 8730
rect 2432 8676 2488 8678
rect 2512 8676 2568 8678
rect 2592 8676 2648 8678
rect 2672 8676 2728 8678
rect 4065 8730 4121 8732
rect 4145 8730 4201 8732
rect 4225 8730 4281 8732
rect 4305 8730 4361 8732
rect 4065 8678 4111 8730
rect 4111 8678 4121 8730
rect 4145 8678 4175 8730
rect 4175 8678 4187 8730
rect 4187 8678 4201 8730
rect 4225 8678 4239 8730
rect 4239 8678 4251 8730
rect 4251 8678 4281 8730
rect 4305 8678 4315 8730
rect 4315 8678 4361 8730
rect 4065 8676 4121 8678
rect 4145 8676 4201 8678
rect 4225 8676 4281 8678
rect 4305 8676 4361 8678
rect 5698 8730 5754 8732
rect 5778 8730 5834 8732
rect 5858 8730 5914 8732
rect 5938 8730 5994 8732
rect 5698 8678 5744 8730
rect 5744 8678 5754 8730
rect 5778 8678 5808 8730
rect 5808 8678 5820 8730
rect 5820 8678 5834 8730
rect 5858 8678 5872 8730
rect 5872 8678 5884 8730
rect 5884 8678 5914 8730
rect 5938 8678 5948 8730
rect 5948 8678 5994 8730
rect 5698 8676 5754 8678
rect 5778 8676 5834 8678
rect 5858 8676 5914 8678
rect 5938 8676 5994 8678
rect 7331 8730 7387 8732
rect 7411 8730 7467 8732
rect 7491 8730 7547 8732
rect 7571 8730 7627 8732
rect 7331 8678 7377 8730
rect 7377 8678 7387 8730
rect 7411 8678 7441 8730
rect 7441 8678 7453 8730
rect 7453 8678 7467 8730
rect 7491 8678 7505 8730
rect 7505 8678 7517 8730
rect 7517 8678 7547 8730
rect 7571 8678 7581 8730
rect 7581 8678 7627 8730
rect 7331 8676 7387 8678
rect 7411 8676 7467 8678
rect 7491 8676 7547 8678
rect 7571 8676 7627 8678
rect 1772 8186 1828 8188
rect 1852 8186 1908 8188
rect 1932 8186 1988 8188
rect 2012 8186 2068 8188
rect 1772 8134 1818 8186
rect 1818 8134 1828 8186
rect 1852 8134 1882 8186
rect 1882 8134 1894 8186
rect 1894 8134 1908 8186
rect 1932 8134 1946 8186
rect 1946 8134 1958 8186
rect 1958 8134 1988 8186
rect 2012 8134 2022 8186
rect 2022 8134 2068 8186
rect 1772 8132 1828 8134
rect 1852 8132 1908 8134
rect 1932 8132 1988 8134
rect 2012 8132 2068 8134
rect 3405 8186 3461 8188
rect 3485 8186 3541 8188
rect 3565 8186 3621 8188
rect 3645 8186 3701 8188
rect 3405 8134 3451 8186
rect 3451 8134 3461 8186
rect 3485 8134 3515 8186
rect 3515 8134 3527 8186
rect 3527 8134 3541 8186
rect 3565 8134 3579 8186
rect 3579 8134 3591 8186
rect 3591 8134 3621 8186
rect 3645 8134 3655 8186
rect 3655 8134 3701 8186
rect 3405 8132 3461 8134
rect 3485 8132 3541 8134
rect 3565 8132 3621 8134
rect 3645 8132 3701 8134
rect 2432 7642 2488 7644
rect 2512 7642 2568 7644
rect 2592 7642 2648 7644
rect 2672 7642 2728 7644
rect 2432 7590 2478 7642
rect 2478 7590 2488 7642
rect 2512 7590 2542 7642
rect 2542 7590 2554 7642
rect 2554 7590 2568 7642
rect 2592 7590 2606 7642
rect 2606 7590 2618 7642
rect 2618 7590 2648 7642
rect 2672 7590 2682 7642
rect 2682 7590 2728 7642
rect 2432 7588 2488 7590
rect 2512 7588 2568 7590
rect 2592 7588 2648 7590
rect 2672 7588 2728 7590
rect 4065 7642 4121 7644
rect 4145 7642 4201 7644
rect 4225 7642 4281 7644
rect 4305 7642 4361 7644
rect 4065 7590 4111 7642
rect 4111 7590 4121 7642
rect 4145 7590 4175 7642
rect 4175 7590 4187 7642
rect 4187 7590 4201 7642
rect 4225 7590 4239 7642
rect 4239 7590 4251 7642
rect 4251 7590 4281 7642
rect 4305 7590 4315 7642
rect 4315 7590 4361 7642
rect 4065 7588 4121 7590
rect 4145 7588 4201 7590
rect 4225 7588 4281 7590
rect 4305 7588 4361 7590
rect 1772 7098 1828 7100
rect 1852 7098 1908 7100
rect 1932 7098 1988 7100
rect 2012 7098 2068 7100
rect 1772 7046 1818 7098
rect 1818 7046 1828 7098
rect 1852 7046 1882 7098
rect 1882 7046 1894 7098
rect 1894 7046 1908 7098
rect 1932 7046 1946 7098
rect 1946 7046 1958 7098
rect 1958 7046 1988 7098
rect 2012 7046 2022 7098
rect 2022 7046 2068 7098
rect 1772 7044 1828 7046
rect 1852 7044 1908 7046
rect 1932 7044 1988 7046
rect 2012 7044 2068 7046
rect 1398 6840 1454 6896
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 1772 6010 1828 6012
rect 1852 6010 1908 6012
rect 1932 6010 1988 6012
rect 2012 6010 2068 6012
rect 1772 5958 1818 6010
rect 1818 5958 1828 6010
rect 1852 5958 1882 6010
rect 1882 5958 1894 6010
rect 1894 5958 1908 6010
rect 1932 5958 1946 6010
rect 1946 5958 1958 6010
rect 1958 5958 1988 6010
rect 2012 5958 2022 6010
rect 2022 5958 2068 6010
rect 1772 5956 1828 5958
rect 1852 5956 1908 5958
rect 1932 5956 1988 5958
rect 2012 5956 2068 5958
rect 2432 6554 2488 6556
rect 2512 6554 2568 6556
rect 2592 6554 2648 6556
rect 2672 6554 2728 6556
rect 2432 6502 2478 6554
rect 2478 6502 2488 6554
rect 2512 6502 2542 6554
rect 2542 6502 2554 6554
rect 2554 6502 2568 6554
rect 2592 6502 2606 6554
rect 2606 6502 2618 6554
rect 2618 6502 2648 6554
rect 2672 6502 2682 6554
rect 2682 6502 2728 6554
rect 2432 6500 2488 6502
rect 2512 6500 2568 6502
rect 2592 6500 2648 6502
rect 2672 6500 2728 6502
rect 2432 5466 2488 5468
rect 2512 5466 2568 5468
rect 2592 5466 2648 5468
rect 2672 5466 2728 5468
rect 2432 5414 2478 5466
rect 2478 5414 2488 5466
rect 2512 5414 2542 5466
rect 2542 5414 2554 5466
rect 2554 5414 2568 5466
rect 2592 5414 2606 5466
rect 2606 5414 2618 5466
rect 2618 5414 2648 5466
rect 2672 5414 2682 5466
rect 2682 5414 2728 5466
rect 2432 5412 2488 5414
rect 2512 5412 2568 5414
rect 2592 5412 2648 5414
rect 2672 5412 2728 5414
rect 1772 4922 1828 4924
rect 1852 4922 1908 4924
rect 1932 4922 1988 4924
rect 2012 4922 2068 4924
rect 1772 4870 1818 4922
rect 1818 4870 1828 4922
rect 1852 4870 1882 4922
rect 1882 4870 1894 4922
rect 1894 4870 1908 4922
rect 1932 4870 1946 4922
rect 1946 4870 1958 4922
rect 1958 4870 1988 4922
rect 2012 4870 2022 4922
rect 2022 4870 2068 4922
rect 1772 4868 1828 4870
rect 1852 4868 1908 4870
rect 1932 4868 1988 4870
rect 2012 4868 2068 4870
rect 2432 4378 2488 4380
rect 2512 4378 2568 4380
rect 2592 4378 2648 4380
rect 2672 4378 2728 4380
rect 2432 4326 2478 4378
rect 2478 4326 2488 4378
rect 2512 4326 2542 4378
rect 2542 4326 2554 4378
rect 2554 4326 2568 4378
rect 2592 4326 2606 4378
rect 2606 4326 2618 4378
rect 2618 4326 2648 4378
rect 2672 4326 2682 4378
rect 2682 4326 2728 4378
rect 2432 4324 2488 4326
rect 2512 4324 2568 4326
rect 2592 4324 2648 4326
rect 2672 4324 2728 4326
rect 1772 3834 1828 3836
rect 1852 3834 1908 3836
rect 1932 3834 1988 3836
rect 2012 3834 2068 3836
rect 1772 3782 1818 3834
rect 1818 3782 1828 3834
rect 1852 3782 1882 3834
rect 1882 3782 1894 3834
rect 1894 3782 1908 3834
rect 1932 3782 1946 3834
rect 1946 3782 1958 3834
rect 1958 3782 1988 3834
rect 2012 3782 2022 3834
rect 2022 3782 2068 3834
rect 1772 3780 1828 3782
rect 1852 3780 1908 3782
rect 1932 3780 1988 3782
rect 2012 3780 2068 3782
rect 2432 3290 2488 3292
rect 2512 3290 2568 3292
rect 2592 3290 2648 3292
rect 2672 3290 2728 3292
rect 2432 3238 2478 3290
rect 2478 3238 2488 3290
rect 2512 3238 2542 3290
rect 2542 3238 2554 3290
rect 2554 3238 2568 3290
rect 2592 3238 2606 3290
rect 2606 3238 2618 3290
rect 2618 3238 2648 3290
rect 2672 3238 2682 3290
rect 2682 3238 2728 3290
rect 2432 3236 2488 3238
rect 2512 3236 2568 3238
rect 2592 3236 2648 3238
rect 2672 3236 2728 3238
rect 3405 7098 3461 7100
rect 3485 7098 3541 7100
rect 3565 7098 3621 7100
rect 3645 7098 3701 7100
rect 3405 7046 3451 7098
rect 3451 7046 3461 7098
rect 3485 7046 3515 7098
rect 3515 7046 3527 7098
rect 3527 7046 3541 7098
rect 3565 7046 3579 7098
rect 3579 7046 3591 7098
rect 3591 7046 3621 7098
rect 3645 7046 3655 7098
rect 3655 7046 3701 7098
rect 3405 7044 3461 7046
rect 3485 7044 3541 7046
rect 3565 7044 3621 7046
rect 3645 7044 3701 7046
rect 5038 8186 5094 8188
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5038 8134 5084 8186
rect 5084 8134 5094 8186
rect 5118 8134 5148 8186
rect 5148 8134 5160 8186
rect 5160 8134 5174 8186
rect 5198 8134 5212 8186
rect 5212 8134 5224 8186
rect 5224 8134 5254 8186
rect 5278 8134 5288 8186
rect 5288 8134 5334 8186
rect 5038 8132 5094 8134
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 6671 8186 6727 8188
rect 6751 8186 6807 8188
rect 6831 8186 6887 8188
rect 6911 8186 6967 8188
rect 6671 8134 6717 8186
rect 6717 8134 6727 8186
rect 6751 8134 6781 8186
rect 6781 8134 6793 8186
rect 6793 8134 6807 8186
rect 6831 8134 6845 8186
rect 6845 8134 6857 8186
rect 6857 8134 6887 8186
rect 6911 8134 6921 8186
rect 6921 8134 6967 8186
rect 6671 8132 6727 8134
rect 6751 8132 6807 8134
rect 6831 8132 6887 8134
rect 6911 8132 6967 8134
rect 5698 7642 5754 7644
rect 5778 7642 5834 7644
rect 5858 7642 5914 7644
rect 5938 7642 5994 7644
rect 5698 7590 5744 7642
rect 5744 7590 5754 7642
rect 5778 7590 5808 7642
rect 5808 7590 5820 7642
rect 5820 7590 5834 7642
rect 5858 7590 5872 7642
rect 5872 7590 5884 7642
rect 5884 7590 5914 7642
rect 5938 7590 5948 7642
rect 5948 7590 5994 7642
rect 5698 7588 5754 7590
rect 5778 7588 5834 7590
rect 5858 7588 5914 7590
rect 5938 7588 5994 7590
rect 5038 7098 5094 7100
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5038 7046 5084 7098
rect 5084 7046 5094 7098
rect 5118 7046 5148 7098
rect 5148 7046 5160 7098
rect 5160 7046 5174 7098
rect 5198 7046 5212 7098
rect 5212 7046 5224 7098
rect 5224 7046 5254 7098
rect 5278 7046 5288 7098
rect 5288 7046 5334 7098
rect 5038 7044 5094 7046
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 4618 6740 4620 6760
rect 4620 6740 4672 6760
rect 4672 6740 4674 6760
rect 4618 6704 4674 6740
rect 4065 6554 4121 6556
rect 4145 6554 4201 6556
rect 4225 6554 4281 6556
rect 4305 6554 4361 6556
rect 4065 6502 4111 6554
rect 4111 6502 4121 6554
rect 4145 6502 4175 6554
rect 4175 6502 4187 6554
rect 4187 6502 4201 6554
rect 4225 6502 4239 6554
rect 4239 6502 4251 6554
rect 4251 6502 4281 6554
rect 4305 6502 4315 6554
rect 4315 6502 4361 6554
rect 4065 6500 4121 6502
rect 4145 6500 4201 6502
rect 4225 6500 4281 6502
rect 4305 6500 4361 6502
rect 3405 6010 3461 6012
rect 3485 6010 3541 6012
rect 3565 6010 3621 6012
rect 3645 6010 3701 6012
rect 3405 5958 3451 6010
rect 3451 5958 3461 6010
rect 3485 5958 3515 6010
rect 3515 5958 3527 6010
rect 3527 5958 3541 6010
rect 3565 5958 3579 6010
rect 3579 5958 3591 6010
rect 3591 5958 3621 6010
rect 3645 5958 3655 6010
rect 3655 5958 3701 6010
rect 3405 5956 3461 5958
rect 3485 5956 3541 5958
rect 3565 5956 3621 5958
rect 3645 5956 3701 5958
rect 4065 5466 4121 5468
rect 4145 5466 4201 5468
rect 4225 5466 4281 5468
rect 4305 5466 4361 5468
rect 4065 5414 4111 5466
rect 4111 5414 4121 5466
rect 4145 5414 4175 5466
rect 4175 5414 4187 5466
rect 4187 5414 4201 5466
rect 4225 5414 4239 5466
rect 4239 5414 4251 5466
rect 4251 5414 4281 5466
rect 4305 5414 4315 5466
rect 4315 5414 4361 5466
rect 4065 5412 4121 5414
rect 4145 5412 4201 5414
rect 4225 5412 4281 5414
rect 4305 5412 4361 5414
rect 7331 7642 7387 7644
rect 7411 7642 7467 7644
rect 7491 7642 7547 7644
rect 7571 7642 7627 7644
rect 7331 7590 7377 7642
rect 7377 7590 7387 7642
rect 7411 7590 7441 7642
rect 7441 7590 7453 7642
rect 7453 7590 7467 7642
rect 7491 7590 7505 7642
rect 7505 7590 7517 7642
rect 7517 7590 7547 7642
rect 7571 7590 7581 7642
rect 7581 7590 7627 7642
rect 7331 7588 7387 7590
rect 7411 7588 7467 7590
rect 7491 7588 7547 7590
rect 7571 7588 7627 7590
rect 7746 7520 7802 7576
rect 5630 6740 5632 6760
rect 5632 6740 5684 6760
rect 5684 6740 5686 6760
rect 5630 6704 5686 6740
rect 3405 4922 3461 4924
rect 3485 4922 3541 4924
rect 3565 4922 3621 4924
rect 3645 4922 3701 4924
rect 3405 4870 3451 4922
rect 3451 4870 3461 4922
rect 3485 4870 3515 4922
rect 3515 4870 3527 4922
rect 3527 4870 3541 4922
rect 3565 4870 3579 4922
rect 3579 4870 3591 4922
rect 3591 4870 3621 4922
rect 3645 4870 3655 4922
rect 3655 4870 3701 4922
rect 3405 4868 3461 4870
rect 3485 4868 3541 4870
rect 3565 4868 3621 4870
rect 3645 4868 3701 4870
rect 3405 3834 3461 3836
rect 3485 3834 3541 3836
rect 3565 3834 3621 3836
rect 3645 3834 3701 3836
rect 3405 3782 3451 3834
rect 3451 3782 3461 3834
rect 3485 3782 3515 3834
rect 3515 3782 3527 3834
rect 3527 3782 3541 3834
rect 3565 3782 3579 3834
rect 3579 3782 3591 3834
rect 3591 3782 3621 3834
rect 3645 3782 3655 3834
rect 3655 3782 3701 3834
rect 3405 3780 3461 3782
rect 3485 3780 3541 3782
rect 3565 3780 3621 3782
rect 3645 3780 3701 3782
rect 4065 4378 4121 4380
rect 4145 4378 4201 4380
rect 4225 4378 4281 4380
rect 4305 4378 4361 4380
rect 4065 4326 4111 4378
rect 4111 4326 4121 4378
rect 4145 4326 4175 4378
rect 4175 4326 4187 4378
rect 4187 4326 4201 4378
rect 4225 4326 4239 4378
rect 4239 4326 4251 4378
rect 4251 4326 4281 4378
rect 4305 4326 4315 4378
rect 4315 4326 4361 4378
rect 4065 4324 4121 4326
rect 4145 4324 4201 4326
rect 4225 4324 4281 4326
rect 4305 4324 4361 4326
rect 5038 6010 5094 6012
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5038 5958 5084 6010
rect 5084 5958 5094 6010
rect 5118 5958 5148 6010
rect 5148 5958 5160 6010
rect 5160 5958 5174 6010
rect 5198 5958 5212 6010
rect 5212 5958 5224 6010
rect 5224 5958 5254 6010
rect 5278 5958 5288 6010
rect 5288 5958 5334 6010
rect 5038 5956 5094 5958
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5038 4922 5094 4924
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5038 4870 5084 4922
rect 5084 4870 5094 4922
rect 5118 4870 5148 4922
rect 5148 4870 5160 4922
rect 5160 4870 5174 4922
rect 5198 4870 5212 4922
rect 5212 4870 5224 4922
rect 5224 4870 5254 4922
rect 5278 4870 5288 4922
rect 5288 4870 5334 4922
rect 5038 4868 5094 4870
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5038 3834 5094 3836
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5038 3782 5084 3834
rect 5084 3782 5094 3834
rect 5118 3782 5148 3834
rect 5148 3782 5160 3834
rect 5160 3782 5174 3834
rect 5198 3782 5212 3834
rect 5212 3782 5224 3834
rect 5224 3782 5254 3834
rect 5278 3782 5288 3834
rect 5288 3782 5334 3834
rect 5038 3780 5094 3782
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5698 6554 5754 6556
rect 5778 6554 5834 6556
rect 5858 6554 5914 6556
rect 5938 6554 5994 6556
rect 5698 6502 5744 6554
rect 5744 6502 5754 6554
rect 5778 6502 5808 6554
rect 5808 6502 5820 6554
rect 5820 6502 5834 6554
rect 5858 6502 5872 6554
rect 5872 6502 5884 6554
rect 5884 6502 5914 6554
rect 5938 6502 5948 6554
rect 5948 6502 5994 6554
rect 5698 6500 5754 6502
rect 5778 6500 5834 6502
rect 5858 6500 5914 6502
rect 5938 6500 5994 6502
rect 6671 7098 6727 7100
rect 6751 7098 6807 7100
rect 6831 7098 6887 7100
rect 6911 7098 6967 7100
rect 6671 7046 6717 7098
rect 6717 7046 6727 7098
rect 6751 7046 6781 7098
rect 6781 7046 6793 7098
rect 6793 7046 6807 7098
rect 6831 7046 6845 7098
rect 6845 7046 6857 7098
rect 6857 7046 6887 7098
rect 6911 7046 6921 7098
rect 6921 7046 6967 7098
rect 6671 7044 6727 7046
rect 6751 7044 6807 7046
rect 6831 7044 6887 7046
rect 6911 7044 6967 7046
rect 7194 6840 7250 6896
rect 5722 6316 5778 6352
rect 5722 6296 5724 6316
rect 5724 6296 5776 6316
rect 5776 6296 5778 6316
rect 5698 5466 5754 5468
rect 5778 5466 5834 5468
rect 5858 5466 5914 5468
rect 5938 5466 5994 5468
rect 5698 5414 5744 5466
rect 5744 5414 5754 5466
rect 5778 5414 5808 5466
rect 5808 5414 5820 5466
rect 5820 5414 5834 5466
rect 5858 5414 5872 5466
rect 5872 5414 5884 5466
rect 5884 5414 5914 5466
rect 5938 5414 5948 5466
rect 5948 5414 5994 5466
rect 5698 5412 5754 5414
rect 5778 5412 5834 5414
rect 5858 5412 5914 5414
rect 5938 5412 5994 5414
rect 7331 6554 7387 6556
rect 7411 6554 7467 6556
rect 7491 6554 7547 6556
rect 7571 6554 7627 6556
rect 7331 6502 7377 6554
rect 7377 6502 7387 6554
rect 7411 6502 7441 6554
rect 7441 6502 7453 6554
rect 7453 6502 7467 6554
rect 7491 6502 7505 6554
rect 7505 6502 7517 6554
rect 7517 6502 7547 6554
rect 7571 6502 7581 6554
rect 7581 6502 7627 6554
rect 7331 6500 7387 6502
rect 7411 6500 7467 6502
rect 7491 6500 7547 6502
rect 7571 6500 7627 6502
rect 6734 6296 6790 6352
rect 7286 6160 7342 6216
rect 6671 6010 6727 6012
rect 6751 6010 6807 6012
rect 6831 6010 6887 6012
rect 6911 6010 6967 6012
rect 6671 5958 6717 6010
rect 6717 5958 6727 6010
rect 6751 5958 6781 6010
rect 6781 5958 6793 6010
rect 6793 5958 6807 6010
rect 6831 5958 6845 6010
rect 6845 5958 6857 6010
rect 6857 5958 6887 6010
rect 6911 5958 6921 6010
rect 6921 5958 6967 6010
rect 6671 5956 6727 5958
rect 6751 5956 6807 5958
rect 6831 5956 6887 5958
rect 6911 5956 6967 5958
rect 7746 5480 7802 5536
rect 7331 5466 7387 5468
rect 7411 5466 7467 5468
rect 7491 5466 7547 5468
rect 7571 5466 7627 5468
rect 7331 5414 7377 5466
rect 7377 5414 7387 5466
rect 7411 5414 7441 5466
rect 7441 5414 7453 5466
rect 7453 5414 7467 5466
rect 7491 5414 7505 5466
rect 7505 5414 7517 5466
rect 7517 5414 7547 5466
rect 7571 5414 7581 5466
rect 7581 5414 7627 5466
rect 7331 5412 7387 5414
rect 7411 5412 7467 5414
rect 7491 5412 7547 5414
rect 7571 5412 7627 5414
rect 6671 4922 6727 4924
rect 6751 4922 6807 4924
rect 6831 4922 6887 4924
rect 6911 4922 6967 4924
rect 6671 4870 6717 4922
rect 6717 4870 6727 4922
rect 6751 4870 6781 4922
rect 6781 4870 6793 4922
rect 6793 4870 6807 4922
rect 6831 4870 6845 4922
rect 6845 4870 6857 4922
rect 6857 4870 6887 4922
rect 6911 4870 6921 4922
rect 6921 4870 6967 4922
rect 6671 4868 6727 4870
rect 6751 4868 6807 4870
rect 6831 4868 6887 4870
rect 6911 4868 6967 4870
rect 7194 4800 7250 4856
rect 5698 4378 5754 4380
rect 5778 4378 5834 4380
rect 5858 4378 5914 4380
rect 5938 4378 5994 4380
rect 5698 4326 5744 4378
rect 5744 4326 5754 4378
rect 5778 4326 5808 4378
rect 5808 4326 5820 4378
rect 5820 4326 5834 4378
rect 5858 4326 5872 4378
rect 5872 4326 5884 4378
rect 5884 4326 5914 4378
rect 5938 4326 5948 4378
rect 5948 4326 5994 4378
rect 5698 4324 5754 4326
rect 5778 4324 5834 4326
rect 5858 4324 5914 4326
rect 5938 4324 5994 4326
rect 7331 4378 7387 4380
rect 7411 4378 7467 4380
rect 7491 4378 7547 4380
rect 7571 4378 7627 4380
rect 7331 4326 7377 4378
rect 7377 4326 7387 4378
rect 7411 4326 7441 4378
rect 7441 4326 7453 4378
rect 7453 4326 7467 4378
rect 7491 4326 7505 4378
rect 7505 4326 7517 4378
rect 7517 4326 7547 4378
rect 7571 4326 7581 4378
rect 7581 4326 7627 4378
rect 7331 4324 7387 4326
rect 7411 4324 7467 4326
rect 7491 4324 7547 4326
rect 7571 4324 7627 4326
rect 7746 4120 7802 4176
rect 6671 3834 6727 3836
rect 6751 3834 6807 3836
rect 6831 3834 6887 3836
rect 6911 3834 6967 3836
rect 6671 3782 6717 3834
rect 6717 3782 6727 3834
rect 6751 3782 6781 3834
rect 6781 3782 6793 3834
rect 6793 3782 6807 3834
rect 6831 3782 6845 3834
rect 6845 3782 6857 3834
rect 6857 3782 6887 3834
rect 6911 3782 6921 3834
rect 6921 3782 6967 3834
rect 6671 3780 6727 3782
rect 6751 3780 6807 3782
rect 6831 3780 6887 3782
rect 6911 3780 6967 3782
rect 4065 3290 4121 3292
rect 4145 3290 4201 3292
rect 4225 3290 4281 3292
rect 4305 3290 4361 3292
rect 4065 3238 4111 3290
rect 4111 3238 4121 3290
rect 4145 3238 4175 3290
rect 4175 3238 4187 3290
rect 4187 3238 4201 3290
rect 4225 3238 4239 3290
rect 4239 3238 4251 3290
rect 4251 3238 4281 3290
rect 4305 3238 4315 3290
rect 4315 3238 4361 3290
rect 4065 3236 4121 3238
rect 4145 3236 4201 3238
rect 4225 3236 4281 3238
rect 4305 3236 4361 3238
rect 1772 2746 1828 2748
rect 1852 2746 1908 2748
rect 1932 2746 1988 2748
rect 2012 2746 2068 2748
rect 1772 2694 1818 2746
rect 1818 2694 1828 2746
rect 1852 2694 1882 2746
rect 1882 2694 1894 2746
rect 1894 2694 1908 2746
rect 1932 2694 1946 2746
rect 1946 2694 1958 2746
rect 1958 2694 1988 2746
rect 2012 2694 2022 2746
rect 2022 2694 2068 2746
rect 1772 2692 1828 2694
rect 1852 2692 1908 2694
rect 1932 2692 1988 2694
rect 2012 2692 2068 2694
rect 3405 2746 3461 2748
rect 3485 2746 3541 2748
rect 3565 2746 3621 2748
rect 3645 2746 3701 2748
rect 3405 2694 3451 2746
rect 3451 2694 3461 2746
rect 3485 2694 3515 2746
rect 3515 2694 3527 2746
rect 3527 2694 3541 2746
rect 3565 2694 3579 2746
rect 3579 2694 3591 2746
rect 3591 2694 3621 2746
rect 3645 2694 3655 2746
rect 3655 2694 3701 2746
rect 3405 2692 3461 2694
rect 3485 2692 3541 2694
rect 3565 2692 3621 2694
rect 3645 2692 3701 2694
rect 5698 3290 5754 3292
rect 5778 3290 5834 3292
rect 5858 3290 5914 3292
rect 5938 3290 5994 3292
rect 5698 3238 5744 3290
rect 5744 3238 5754 3290
rect 5778 3238 5808 3290
rect 5808 3238 5820 3290
rect 5820 3238 5834 3290
rect 5858 3238 5872 3290
rect 5872 3238 5884 3290
rect 5884 3238 5914 3290
rect 5938 3238 5948 3290
rect 5948 3238 5994 3290
rect 5698 3236 5754 3238
rect 5778 3236 5834 3238
rect 5858 3236 5914 3238
rect 5938 3236 5994 3238
rect 7194 3440 7250 3496
rect 7331 3290 7387 3292
rect 7411 3290 7467 3292
rect 7491 3290 7547 3292
rect 7571 3290 7627 3292
rect 7331 3238 7377 3290
rect 7377 3238 7387 3290
rect 7411 3238 7441 3290
rect 7441 3238 7453 3290
rect 7453 3238 7467 3290
rect 7491 3238 7505 3290
rect 7505 3238 7517 3290
rect 7517 3238 7547 3290
rect 7571 3238 7581 3290
rect 7581 3238 7627 3290
rect 7331 3236 7387 3238
rect 7411 3236 7467 3238
rect 7491 3236 7547 3238
rect 7571 3236 7627 3238
rect 7286 2760 7342 2816
rect 5038 2746 5094 2748
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5038 2694 5084 2746
rect 5084 2694 5094 2746
rect 5118 2694 5148 2746
rect 5148 2694 5160 2746
rect 5160 2694 5174 2746
rect 5198 2694 5212 2746
rect 5212 2694 5224 2746
rect 5224 2694 5254 2746
rect 5278 2694 5288 2746
rect 5288 2694 5334 2746
rect 5038 2692 5094 2694
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 6671 2746 6727 2748
rect 6751 2746 6807 2748
rect 6831 2746 6887 2748
rect 6911 2746 6967 2748
rect 6671 2694 6717 2746
rect 6717 2694 6727 2746
rect 6751 2694 6781 2746
rect 6781 2694 6793 2746
rect 6793 2694 6807 2746
rect 6831 2694 6845 2746
rect 6845 2694 6857 2746
rect 6857 2694 6887 2746
rect 6911 2694 6921 2746
rect 6921 2694 6967 2746
rect 6671 2692 6727 2694
rect 6751 2692 6807 2694
rect 6831 2692 6887 2694
rect 6911 2692 6967 2694
rect 2432 2202 2488 2204
rect 2512 2202 2568 2204
rect 2592 2202 2648 2204
rect 2672 2202 2728 2204
rect 2432 2150 2478 2202
rect 2478 2150 2488 2202
rect 2512 2150 2542 2202
rect 2542 2150 2554 2202
rect 2554 2150 2568 2202
rect 2592 2150 2606 2202
rect 2606 2150 2618 2202
rect 2618 2150 2648 2202
rect 2672 2150 2682 2202
rect 2682 2150 2728 2202
rect 2432 2148 2488 2150
rect 2512 2148 2568 2150
rect 2592 2148 2648 2150
rect 2672 2148 2728 2150
rect 4065 2202 4121 2204
rect 4145 2202 4201 2204
rect 4225 2202 4281 2204
rect 4305 2202 4361 2204
rect 4065 2150 4111 2202
rect 4111 2150 4121 2202
rect 4145 2150 4175 2202
rect 4175 2150 4187 2202
rect 4187 2150 4201 2202
rect 4225 2150 4239 2202
rect 4239 2150 4251 2202
rect 4251 2150 4281 2202
rect 4305 2150 4315 2202
rect 4315 2150 4361 2202
rect 4065 2148 4121 2150
rect 4145 2148 4201 2150
rect 4225 2148 4281 2150
rect 4305 2148 4361 2150
rect 5698 2202 5754 2204
rect 5778 2202 5834 2204
rect 5858 2202 5914 2204
rect 5938 2202 5994 2204
rect 5698 2150 5744 2202
rect 5744 2150 5754 2202
rect 5778 2150 5808 2202
rect 5808 2150 5820 2202
rect 5820 2150 5834 2202
rect 5858 2150 5872 2202
rect 5872 2150 5884 2202
rect 5884 2150 5914 2202
rect 5938 2150 5948 2202
rect 5948 2150 5994 2202
rect 5698 2148 5754 2150
rect 5778 2148 5834 2150
rect 5858 2148 5914 2150
rect 5938 2148 5994 2150
rect 7331 2202 7387 2204
rect 7411 2202 7467 2204
rect 7491 2202 7547 2204
rect 7571 2202 7627 2204
rect 7331 2150 7377 2202
rect 7377 2150 7387 2202
rect 7411 2150 7441 2202
rect 7441 2150 7453 2202
rect 7453 2150 7467 2202
rect 7491 2150 7505 2202
rect 7505 2150 7517 2202
rect 7517 2150 7547 2202
rect 7571 2150 7581 2202
rect 7581 2150 7627 2202
rect 7331 2148 7387 2150
rect 7411 2148 7467 2150
rect 7491 2148 7547 2150
rect 7571 2148 7627 2150
<< metal3 >>
rect 2422 8736 2738 8737
rect 2422 8672 2428 8736
rect 2492 8672 2508 8736
rect 2572 8672 2588 8736
rect 2652 8672 2668 8736
rect 2732 8672 2738 8736
rect 2422 8671 2738 8672
rect 4055 8736 4371 8737
rect 4055 8672 4061 8736
rect 4125 8672 4141 8736
rect 4205 8672 4221 8736
rect 4285 8672 4301 8736
rect 4365 8672 4371 8736
rect 4055 8671 4371 8672
rect 5688 8736 6004 8737
rect 5688 8672 5694 8736
rect 5758 8672 5774 8736
rect 5838 8672 5854 8736
rect 5918 8672 5934 8736
rect 5998 8672 6004 8736
rect 5688 8671 6004 8672
rect 7321 8736 7637 8737
rect 7321 8672 7327 8736
rect 7391 8672 7407 8736
rect 7471 8672 7487 8736
rect 7551 8672 7567 8736
rect 7631 8672 7637 8736
rect 7321 8671 7637 8672
rect 1762 8192 2078 8193
rect 1762 8128 1768 8192
rect 1832 8128 1848 8192
rect 1912 8128 1928 8192
rect 1992 8128 2008 8192
rect 2072 8128 2078 8192
rect 1762 8127 2078 8128
rect 3395 8192 3711 8193
rect 3395 8128 3401 8192
rect 3465 8128 3481 8192
rect 3545 8128 3561 8192
rect 3625 8128 3641 8192
rect 3705 8128 3711 8192
rect 3395 8127 3711 8128
rect 5028 8192 5344 8193
rect 5028 8128 5034 8192
rect 5098 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5344 8192
rect 5028 8127 5344 8128
rect 6661 8192 6977 8193
rect 6661 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6907 8192
rect 6971 8128 6977 8192
rect 6661 8127 6977 8128
rect 2422 7648 2738 7649
rect 2422 7584 2428 7648
rect 2492 7584 2508 7648
rect 2572 7584 2588 7648
rect 2652 7584 2668 7648
rect 2732 7584 2738 7648
rect 2422 7583 2738 7584
rect 4055 7648 4371 7649
rect 4055 7584 4061 7648
rect 4125 7584 4141 7648
rect 4205 7584 4221 7648
rect 4285 7584 4301 7648
rect 4365 7584 4371 7648
rect 4055 7583 4371 7584
rect 5688 7648 6004 7649
rect 5688 7584 5694 7648
rect 5758 7584 5774 7648
rect 5838 7584 5854 7648
rect 5918 7584 5934 7648
rect 5998 7584 6004 7648
rect 5688 7583 6004 7584
rect 7321 7648 7637 7649
rect 7321 7584 7327 7648
rect 7391 7584 7407 7648
rect 7471 7584 7487 7648
rect 7551 7584 7567 7648
rect 7631 7584 7637 7648
rect 7321 7583 7637 7584
rect 7741 7578 7807 7581
rect 8019 7578 8819 7608
rect 7741 7576 8819 7578
rect 7741 7520 7746 7576
rect 7802 7520 8819 7576
rect 7741 7518 8819 7520
rect 7741 7515 7807 7518
rect 8019 7488 8819 7518
rect 1762 7104 2078 7105
rect 1762 7040 1768 7104
rect 1832 7040 1848 7104
rect 1912 7040 1928 7104
rect 1992 7040 2008 7104
rect 2072 7040 2078 7104
rect 1762 7039 2078 7040
rect 3395 7104 3711 7105
rect 3395 7040 3401 7104
rect 3465 7040 3481 7104
rect 3545 7040 3561 7104
rect 3625 7040 3641 7104
rect 3705 7040 3711 7104
rect 3395 7039 3711 7040
rect 5028 7104 5344 7105
rect 5028 7040 5034 7104
rect 5098 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5344 7104
rect 5028 7039 5344 7040
rect 6661 7104 6977 7105
rect 6661 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6907 7104
rect 6971 7040 6977 7104
rect 6661 7039 6977 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 7189 6898 7255 6901
rect 8019 6898 8819 6928
rect 7189 6896 8819 6898
rect 7189 6840 7194 6896
rect 7250 6840 8819 6896
rect 7189 6838 8819 6840
rect 7189 6835 7255 6838
rect 8019 6808 8819 6838
rect 4613 6762 4679 6765
rect 5625 6762 5691 6765
rect 4613 6760 5691 6762
rect 4613 6704 4618 6760
rect 4674 6704 5630 6760
rect 5686 6704 5691 6760
rect 4613 6702 5691 6704
rect 4613 6699 4679 6702
rect 5625 6699 5691 6702
rect 2422 6560 2738 6561
rect 2422 6496 2428 6560
rect 2492 6496 2508 6560
rect 2572 6496 2588 6560
rect 2652 6496 2668 6560
rect 2732 6496 2738 6560
rect 2422 6495 2738 6496
rect 4055 6560 4371 6561
rect 4055 6496 4061 6560
rect 4125 6496 4141 6560
rect 4205 6496 4221 6560
rect 4285 6496 4301 6560
rect 4365 6496 4371 6560
rect 4055 6495 4371 6496
rect 5688 6560 6004 6561
rect 5688 6496 5694 6560
rect 5758 6496 5774 6560
rect 5838 6496 5854 6560
rect 5918 6496 5934 6560
rect 5998 6496 6004 6560
rect 5688 6495 6004 6496
rect 7321 6560 7637 6561
rect 7321 6496 7327 6560
rect 7391 6496 7407 6560
rect 7471 6496 7487 6560
rect 7551 6496 7567 6560
rect 7631 6496 7637 6560
rect 7321 6495 7637 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 5717 6354 5783 6357
rect 6729 6354 6795 6357
rect 5717 6352 6795 6354
rect 5717 6296 5722 6352
rect 5778 6296 6734 6352
rect 6790 6296 6795 6352
rect 5717 6294 6795 6296
rect 5717 6291 5783 6294
rect 6729 6291 6795 6294
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 7281 6218 7347 6221
rect 8019 6218 8819 6248
rect 7281 6216 8819 6218
rect 7281 6160 7286 6216
rect 7342 6160 8819 6216
rect 7281 6158 8819 6160
rect 0 6128 800 6158
rect 7281 6155 7347 6158
rect 8019 6128 8819 6158
rect 1762 6016 2078 6017
rect 1762 5952 1768 6016
rect 1832 5952 1848 6016
rect 1912 5952 1928 6016
rect 1992 5952 2008 6016
rect 2072 5952 2078 6016
rect 1762 5951 2078 5952
rect 3395 6016 3711 6017
rect 3395 5952 3401 6016
rect 3465 5952 3481 6016
rect 3545 5952 3561 6016
rect 3625 5952 3641 6016
rect 3705 5952 3711 6016
rect 3395 5951 3711 5952
rect 5028 6016 5344 6017
rect 5028 5952 5034 6016
rect 5098 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5344 6016
rect 5028 5951 5344 5952
rect 6661 6016 6977 6017
rect 6661 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6907 6016
rect 6971 5952 6977 6016
rect 6661 5951 6977 5952
rect 7741 5538 7807 5541
rect 8019 5538 8819 5568
rect 7741 5536 8819 5538
rect 7741 5480 7746 5536
rect 7802 5480 8819 5536
rect 7741 5478 8819 5480
rect 7741 5475 7807 5478
rect 2422 5472 2738 5473
rect 2422 5408 2428 5472
rect 2492 5408 2508 5472
rect 2572 5408 2588 5472
rect 2652 5408 2668 5472
rect 2732 5408 2738 5472
rect 2422 5407 2738 5408
rect 4055 5472 4371 5473
rect 4055 5408 4061 5472
rect 4125 5408 4141 5472
rect 4205 5408 4221 5472
rect 4285 5408 4301 5472
rect 4365 5408 4371 5472
rect 4055 5407 4371 5408
rect 5688 5472 6004 5473
rect 5688 5408 5694 5472
rect 5758 5408 5774 5472
rect 5838 5408 5854 5472
rect 5918 5408 5934 5472
rect 5998 5408 6004 5472
rect 5688 5407 6004 5408
rect 7321 5472 7637 5473
rect 7321 5408 7327 5472
rect 7391 5408 7407 5472
rect 7471 5408 7487 5472
rect 7551 5408 7567 5472
rect 7631 5408 7637 5472
rect 8019 5448 8819 5478
rect 7321 5407 7637 5408
rect 1762 4928 2078 4929
rect 1762 4864 1768 4928
rect 1832 4864 1848 4928
rect 1912 4864 1928 4928
rect 1992 4864 2008 4928
rect 2072 4864 2078 4928
rect 1762 4863 2078 4864
rect 3395 4928 3711 4929
rect 3395 4864 3401 4928
rect 3465 4864 3481 4928
rect 3545 4864 3561 4928
rect 3625 4864 3641 4928
rect 3705 4864 3711 4928
rect 3395 4863 3711 4864
rect 5028 4928 5344 4929
rect 5028 4864 5034 4928
rect 5098 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5344 4928
rect 5028 4863 5344 4864
rect 6661 4928 6977 4929
rect 6661 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6907 4928
rect 6971 4864 6977 4928
rect 6661 4863 6977 4864
rect 7189 4858 7255 4861
rect 8019 4858 8819 4888
rect 7189 4856 8819 4858
rect 7189 4800 7194 4856
rect 7250 4800 8819 4856
rect 7189 4798 8819 4800
rect 7189 4795 7255 4798
rect 8019 4768 8819 4798
rect 2422 4384 2738 4385
rect 2422 4320 2428 4384
rect 2492 4320 2508 4384
rect 2572 4320 2588 4384
rect 2652 4320 2668 4384
rect 2732 4320 2738 4384
rect 2422 4319 2738 4320
rect 4055 4384 4371 4385
rect 4055 4320 4061 4384
rect 4125 4320 4141 4384
rect 4205 4320 4221 4384
rect 4285 4320 4301 4384
rect 4365 4320 4371 4384
rect 4055 4319 4371 4320
rect 5688 4384 6004 4385
rect 5688 4320 5694 4384
rect 5758 4320 5774 4384
rect 5838 4320 5854 4384
rect 5918 4320 5934 4384
rect 5998 4320 6004 4384
rect 5688 4319 6004 4320
rect 7321 4384 7637 4385
rect 7321 4320 7327 4384
rect 7391 4320 7407 4384
rect 7471 4320 7487 4384
rect 7551 4320 7567 4384
rect 7631 4320 7637 4384
rect 7321 4319 7637 4320
rect 7741 4178 7807 4181
rect 8019 4178 8819 4208
rect 7741 4176 8819 4178
rect 7741 4120 7746 4176
rect 7802 4120 8819 4176
rect 7741 4118 8819 4120
rect 7741 4115 7807 4118
rect 8019 4088 8819 4118
rect 1762 3840 2078 3841
rect 1762 3776 1768 3840
rect 1832 3776 1848 3840
rect 1912 3776 1928 3840
rect 1992 3776 2008 3840
rect 2072 3776 2078 3840
rect 1762 3775 2078 3776
rect 3395 3840 3711 3841
rect 3395 3776 3401 3840
rect 3465 3776 3481 3840
rect 3545 3776 3561 3840
rect 3625 3776 3641 3840
rect 3705 3776 3711 3840
rect 3395 3775 3711 3776
rect 5028 3840 5344 3841
rect 5028 3776 5034 3840
rect 5098 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5344 3840
rect 5028 3775 5344 3776
rect 6661 3840 6977 3841
rect 6661 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6907 3840
rect 6971 3776 6977 3840
rect 6661 3775 6977 3776
rect 7189 3498 7255 3501
rect 8019 3498 8819 3528
rect 7189 3496 8819 3498
rect 7189 3440 7194 3496
rect 7250 3440 8819 3496
rect 7189 3438 8819 3440
rect 7189 3435 7255 3438
rect 8019 3408 8819 3438
rect 2422 3296 2738 3297
rect 2422 3232 2428 3296
rect 2492 3232 2508 3296
rect 2572 3232 2588 3296
rect 2652 3232 2668 3296
rect 2732 3232 2738 3296
rect 2422 3231 2738 3232
rect 4055 3296 4371 3297
rect 4055 3232 4061 3296
rect 4125 3232 4141 3296
rect 4205 3232 4221 3296
rect 4285 3232 4301 3296
rect 4365 3232 4371 3296
rect 4055 3231 4371 3232
rect 5688 3296 6004 3297
rect 5688 3232 5694 3296
rect 5758 3232 5774 3296
rect 5838 3232 5854 3296
rect 5918 3232 5934 3296
rect 5998 3232 6004 3296
rect 5688 3231 6004 3232
rect 7321 3296 7637 3297
rect 7321 3232 7327 3296
rect 7391 3232 7407 3296
rect 7471 3232 7487 3296
rect 7551 3232 7567 3296
rect 7631 3232 7637 3296
rect 7321 3231 7637 3232
rect 7281 2818 7347 2821
rect 8019 2818 8819 2848
rect 7281 2816 8819 2818
rect 7281 2760 7286 2816
rect 7342 2760 8819 2816
rect 7281 2758 8819 2760
rect 7281 2755 7347 2758
rect 1762 2752 2078 2753
rect 1762 2688 1768 2752
rect 1832 2688 1848 2752
rect 1912 2688 1928 2752
rect 1992 2688 2008 2752
rect 2072 2688 2078 2752
rect 1762 2687 2078 2688
rect 3395 2752 3711 2753
rect 3395 2688 3401 2752
rect 3465 2688 3481 2752
rect 3545 2688 3561 2752
rect 3625 2688 3641 2752
rect 3705 2688 3711 2752
rect 3395 2687 3711 2688
rect 5028 2752 5344 2753
rect 5028 2688 5034 2752
rect 5098 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5344 2752
rect 5028 2687 5344 2688
rect 6661 2752 6977 2753
rect 6661 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6907 2752
rect 6971 2688 6977 2752
rect 8019 2728 8819 2758
rect 6661 2687 6977 2688
rect 2422 2208 2738 2209
rect 2422 2144 2428 2208
rect 2492 2144 2508 2208
rect 2572 2144 2588 2208
rect 2652 2144 2668 2208
rect 2732 2144 2738 2208
rect 2422 2143 2738 2144
rect 4055 2208 4371 2209
rect 4055 2144 4061 2208
rect 4125 2144 4141 2208
rect 4205 2144 4221 2208
rect 4285 2144 4301 2208
rect 4365 2144 4371 2208
rect 4055 2143 4371 2144
rect 5688 2208 6004 2209
rect 5688 2144 5694 2208
rect 5758 2144 5774 2208
rect 5838 2144 5854 2208
rect 5918 2144 5934 2208
rect 5998 2144 6004 2208
rect 5688 2143 6004 2144
rect 7321 2208 7637 2209
rect 7321 2144 7327 2208
rect 7391 2144 7407 2208
rect 7471 2144 7487 2208
rect 7551 2144 7567 2208
rect 7631 2144 7637 2208
rect 7321 2143 7637 2144
<< via3 >>
rect 2428 8732 2492 8736
rect 2428 8676 2432 8732
rect 2432 8676 2488 8732
rect 2488 8676 2492 8732
rect 2428 8672 2492 8676
rect 2508 8732 2572 8736
rect 2508 8676 2512 8732
rect 2512 8676 2568 8732
rect 2568 8676 2572 8732
rect 2508 8672 2572 8676
rect 2588 8732 2652 8736
rect 2588 8676 2592 8732
rect 2592 8676 2648 8732
rect 2648 8676 2652 8732
rect 2588 8672 2652 8676
rect 2668 8732 2732 8736
rect 2668 8676 2672 8732
rect 2672 8676 2728 8732
rect 2728 8676 2732 8732
rect 2668 8672 2732 8676
rect 4061 8732 4125 8736
rect 4061 8676 4065 8732
rect 4065 8676 4121 8732
rect 4121 8676 4125 8732
rect 4061 8672 4125 8676
rect 4141 8732 4205 8736
rect 4141 8676 4145 8732
rect 4145 8676 4201 8732
rect 4201 8676 4205 8732
rect 4141 8672 4205 8676
rect 4221 8732 4285 8736
rect 4221 8676 4225 8732
rect 4225 8676 4281 8732
rect 4281 8676 4285 8732
rect 4221 8672 4285 8676
rect 4301 8732 4365 8736
rect 4301 8676 4305 8732
rect 4305 8676 4361 8732
rect 4361 8676 4365 8732
rect 4301 8672 4365 8676
rect 5694 8732 5758 8736
rect 5694 8676 5698 8732
rect 5698 8676 5754 8732
rect 5754 8676 5758 8732
rect 5694 8672 5758 8676
rect 5774 8732 5838 8736
rect 5774 8676 5778 8732
rect 5778 8676 5834 8732
rect 5834 8676 5838 8732
rect 5774 8672 5838 8676
rect 5854 8732 5918 8736
rect 5854 8676 5858 8732
rect 5858 8676 5914 8732
rect 5914 8676 5918 8732
rect 5854 8672 5918 8676
rect 5934 8732 5998 8736
rect 5934 8676 5938 8732
rect 5938 8676 5994 8732
rect 5994 8676 5998 8732
rect 5934 8672 5998 8676
rect 7327 8732 7391 8736
rect 7327 8676 7331 8732
rect 7331 8676 7387 8732
rect 7387 8676 7391 8732
rect 7327 8672 7391 8676
rect 7407 8732 7471 8736
rect 7407 8676 7411 8732
rect 7411 8676 7467 8732
rect 7467 8676 7471 8732
rect 7407 8672 7471 8676
rect 7487 8732 7551 8736
rect 7487 8676 7491 8732
rect 7491 8676 7547 8732
rect 7547 8676 7551 8732
rect 7487 8672 7551 8676
rect 7567 8732 7631 8736
rect 7567 8676 7571 8732
rect 7571 8676 7627 8732
rect 7627 8676 7631 8732
rect 7567 8672 7631 8676
rect 1768 8188 1832 8192
rect 1768 8132 1772 8188
rect 1772 8132 1828 8188
rect 1828 8132 1832 8188
rect 1768 8128 1832 8132
rect 1848 8188 1912 8192
rect 1848 8132 1852 8188
rect 1852 8132 1908 8188
rect 1908 8132 1912 8188
rect 1848 8128 1912 8132
rect 1928 8188 1992 8192
rect 1928 8132 1932 8188
rect 1932 8132 1988 8188
rect 1988 8132 1992 8188
rect 1928 8128 1992 8132
rect 2008 8188 2072 8192
rect 2008 8132 2012 8188
rect 2012 8132 2068 8188
rect 2068 8132 2072 8188
rect 2008 8128 2072 8132
rect 3401 8188 3465 8192
rect 3401 8132 3405 8188
rect 3405 8132 3461 8188
rect 3461 8132 3465 8188
rect 3401 8128 3465 8132
rect 3481 8188 3545 8192
rect 3481 8132 3485 8188
rect 3485 8132 3541 8188
rect 3541 8132 3545 8188
rect 3481 8128 3545 8132
rect 3561 8188 3625 8192
rect 3561 8132 3565 8188
rect 3565 8132 3621 8188
rect 3621 8132 3625 8188
rect 3561 8128 3625 8132
rect 3641 8188 3705 8192
rect 3641 8132 3645 8188
rect 3645 8132 3701 8188
rect 3701 8132 3705 8188
rect 3641 8128 3705 8132
rect 5034 8188 5098 8192
rect 5034 8132 5038 8188
rect 5038 8132 5094 8188
rect 5094 8132 5098 8188
rect 5034 8128 5098 8132
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 6667 8188 6731 8192
rect 6667 8132 6671 8188
rect 6671 8132 6727 8188
rect 6727 8132 6731 8188
rect 6667 8128 6731 8132
rect 6747 8188 6811 8192
rect 6747 8132 6751 8188
rect 6751 8132 6807 8188
rect 6807 8132 6811 8188
rect 6747 8128 6811 8132
rect 6827 8188 6891 8192
rect 6827 8132 6831 8188
rect 6831 8132 6887 8188
rect 6887 8132 6891 8188
rect 6827 8128 6891 8132
rect 6907 8188 6971 8192
rect 6907 8132 6911 8188
rect 6911 8132 6967 8188
rect 6967 8132 6971 8188
rect 6907 8128 6971 8132
rect 2428 7644 2492 7648
rect 2428 7588 2432 7644
rect 2432 7588 2488 7644
rect 2488 7588 2492 7644
rect 2428 7584 2492 7588
rect 2508 7644 2572 7648
rect 2508 7588 2512 7644
rect 2512 7588 2568 7644
rect 2568 7588 2572 7644
rect 2508 7584 2572 7588
rect 2588 7644 2652 7648
rect 2588 7588 2592 7644
rect 2592 7588 2648 7644
rect 2648 7588 2652 7644
rect 2588 7584 2652 7588
rect 2668 7644 2732 7648
rect 2668 7588 2672 7644
rect 2672 7588 2728 7644
rect 2728 7588 2732 7644
rect 2668 7584 2732 7588
rect 4061 7644 4125 7648
rect 4061 7588 4065 7644
rect 4065 7588 4121 7644
rect 4121 7588 4125 7644
rect 4061 7584 4125 7588
rect 4141 7644 4205 7648
rect 4141 7588 4145 7644
rect 4145 7588 4201 7644
rect 4201 7588 4205 7644
rect 4141 7584 4205 7588
rect 4221 7644 4285 7648
rect 4221 7588 4225 7644
rect 4225 7588 4281 7644
rect 4281 7588 4285 7644
rect 4221 7584 4285 7588
rect 4301 7644 4365 7648
rect 4301 7588 4305 7644
rect 4305 7588 4361 7644
rect 4361 7588 4365 7644
rect 4301 7584 4365 7588
rect 5694 7644 5758 7648
rect 5694 7588 5698 7644
rect 5698 7588 5754 7644
rect 5754 7588 5758 7644
rect 5694 7584 5758 7588
rect 5774 7644 5838 7648
rect 5774 7588 5778 7644
rect 5778 7588 5834 7644
rect 5834 7588 5838 7644
rect 5774 7584 5838 7588
rect 5854 7644 5918 7648
rect 5854 7588 5858 7644
rect 5858 7588 5914 7644
rect 5914 7588 5918 7644
rect 5854 7584 5918 7588
rect 5934 7644 5998 7648
rect 5934 7588 5938 7644
rect 5938 7588 5994 7644
rect 5994 7588 5998 7644
rect 5934 7584 5998 7588
rect 7327 7644 7391 7648
rect 7327 7588 7331 7644
rect 7331 7588 7387 7644
rect 7387 7588 7391 7644
rect 7327 7584 7391 7588
rect 7407 7644 7471 7648
rect 7407 7588 7411 7644
rect 7411 7588 7467 7644
rect 7467 7588 7471 7644
rect 7407 7584 7471 7588
rect 7487 7644 7551 7648
rect 7487 7588 7491 7644
rect 7491 7588 7547 7644
rect 7547 7588 7551 7644
rect 7487 7584 7551 7588
rect 7567 7644 7631 7648
rect 7567 7588 7571 7644
rect 7571 7588 7627 7644
rect 7627 7588 7631 7644
rect 7567 7584 7631 7588
rect 1768 7100 1832 7104
rect 1768 7044 1772 7100
rect 1772 7044 1828 7100
rect 1828 7044 1832 7100
rect 1768 7040 1832 7044
rect 1848 7100 1912 7104
rect 1848 7044 1852 7100
rect 1852 7044 1908 7100
rect 1908 7044 1912 7100
rect 1848 7040 1912 7044
rect 1928 7100 1992 7104
rect 1928 7044 1932 7100
rect 1932 7044 1988 7100
rect 1988 7044 1992 7100
rect 1928 7040 1992 7044
rect 2008 7100 2072 7104
rect 2008 7044 2012 7100
rect 2012 7044 2068 7100
rect 2068 7044 2072 7100
rect 2008 7040 2072 7044
rect 3401 7100 3465 7104
rect 3401 7044 3405 7100
rect 3405 7044 3461 7100
rect 3461 7044 3465 7100
rect 3401 7040 3465 7044
rect 3481 7100 3545 7104
rect 3481 7044 3485 7100
rect 3485 7044 3541 7100
rect 3541 7044 3545 7100
rect 3481 7040 3545 7044
rect 3561 7100 3625 7104
rect 3561 7044 3565 7100
rect 3565 7044 3621 7100
rect 3621 7044 3625 7100
rect 3561 7040 3625 7044
rect 3641 7100 3705 7104
rect 3641 7044 3645 7100
rect 3645 7044 3701 7100
rect 3701 7044 3705 7100
rect 3641 7040 3705 7044
rect 5034 7100 5098 7104
rect 5034 7044 5038 7100
rect 5038 7044 5094 7100
rect 5094 7044 5098 7100
rect 5034 7040 5098 7044
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 6667 7100 6731 7104
rect 6667 7044 6671 7100
rect 6671 7044 6727 7100
rect 6727 7044 6731 7100
rect 6667 7040 6731 7044
rect 6747 7100 6811 7104
rect 6747 7044 6751 7100
rect 6751 7044 6807 7100
rect 6807 7044 6811 7100
rect 6747 7040 6811 7044
rect 6827 7100 6891 7104
rect 6827 7044 6831 7100
rect 6831 7044 6887 7100
rect 6887 7044 6891 7100
rect 6827 7040 6891 7044
rect 6907 7100 6971 7104
rect 6907 7044 6911 7100
rect 6911 7044 6967 7100
rect 6967 7044 6971 7100
rect 6907 7040 6971 7044
rect 2428 6556 2492 6560
rect 2428 6500 2432 6556
rect 2432 6500 2488 6556
rect 2488 6500 2492 6556
rect 2428 6496 2492 6500
rect 2508 6556 2572 6560
rect 2508 6500 2512 6556
rect 2512 6500 2568 6556
rect 2568 6500 2572 6556
rect 2508 6496 2572 6500
rect 2588 6556 2652 6560
rect 2588 6500 2592 6556
rect 2592 6500 2648 6556
rect 2648 6500 2652 6556
rect 2588 6496 2652 6500
rect 2668 6556 2732 6560
rect 2668 6500 2672 6556
rect 2672 6500 2728 6556
rect 2728 6500 2732 6556
rect 2668 6496 2732 6500
rect 4061 6556 4125 6560
rect 4061 6500 4065 6556
rect 4065 6500 4121 6556
rect 4121 6500 4125 6556
rect 4061 6496 4125 6500
rect 4141 6556 4205 6560
rect 4141 6500 4145 6556
rect 4145 6500 4201 6556
rect 4201 6500 4205 6556
rect 4141 6496 4205 6500
rect 4221 6556 4285 6560
rect 4221 6500 4225 6556
rect 4225 6500 4281 6556
rect 4281 6500 4285 6556
rect 4221 6496 4285 6500
rect 4301 6556 4365 6560
rect 4301 6500 4305 6556
rect 4305 6500 4361 6556
rect 4361 6500 4365 6556
rect 4301 6496 4365 6500
rect 5694 6556 5758 6560
rect 5694 6500 5698 6556
rect 5698 6500 5754 6556
rect 5754 6500 5758 6556
rect 5694 6496 5758 6500
rect 5774 6556 5838 6560
rect 5774 6500 5778 6556
rect 5778 6500 5834 6556
rect 5834 6500 5838 6556
rect 5774 6496 5838 6500
rect 5854 6556 5918 6560
rect 5854 6500 5858 6556
rect 5858 6500 5914 6556
rect 5914 6500 5918 6556
rect 5854 6496 5918 6500
rect 5934 6556 5998 6560
rect 5934 6500 5938 6556
rect 5938 6500 5994 6556
rect 5994 6500 5998 6556
rect 5934 6496 5998 6500
rect 7327 6556 7391 6560
rect 7327 6500 7331 6556
rect 7331 6500 7387 6556
rect 7387 6500 7391 6556
rect 7327 6496 7391 6500
rect 7407 6556 7471 6560
rect 7407 6500 7411 6556
rect 7411 6500 7467 6556
rect 7467 6500 7471 6556
rect 7407 6496 7471 6500
rect 7487 6556 7551 6560
rect 7487 6500 7491 6556
rect 7491 6500 7547 6556
rect 7547 6500 7551 6556
rect 7487 6496 7551 6500
rect 7567 6556 7631 6560
rect 7567 6500 7571 6556
rect 7571 6500 7627 6556
rect 7627 6500 7631 6556
rect 7567 6496 7631 6500
rect 1768 6012 1832 6016
rect 1768 5956 1772 6012
rect 1772 5956 1828 6012
rect 1828 5956 1832 6012
rect 1768 5952 1832 5956
rect 1848 6012 1912 6016
rect 1848 5956 1852 6012
rect 1852 5956 1908 6012
rect 1908 5956 1912 6012
rect 1848 5952 1912 5956
rect 1928 6012 1992 6016
rect 1928 5956 1932 6012
rect 1932 5956 1988 6012
rect 1988 5956 1992 6012
rect 1928 5952 1992 5956
rect 2008 6012 2072 6016
rect 2008 5956 2012 6012
rect 2012 5956 2068 6012
rect 2068 5956 2072 6012
rect 2008 5952 2072 5956
rect 3401 6012 3465 6016
rect 3401 5956 3405 6012
rect 3405 5956 3461 6012
rect 3461 5956 3465 6012
rect 3401 5952 3465 5956
rect 3481 6012 3545 6016
rect 3481 5956 3485 6012
rect 3485 5956 3541 6012
rect 3541 5956 3545 6012
rect 3481 5952 3545 5956
rect 3561 6012 3625 6016
rect 3561 5956 3565 6012
rect 3565 5956 3621 6012
rect 3621 5956 3625 6012
rect 3561 5952 3625 5956
rect 3641 6012 3705 6016
rect 3641 5956 3645 6012
rect 3645 5956 3701 6012
rect 3701 5956 3705 6012
rect 3641 5952 3705 5956
rect 5034 6012 5098 6016
rect 5034 5956 5038 6012
rect 5038 5956 5094 6012
rect 5094 5956 5098 6012
rect 5034 5952 5098 5956
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 6667 6012 6731 6016
rect 6667 5956 6671 6012
rect 6671 5956 6727 6012
rect 6727 5956 6731 6012
rect 6667 5952 6731 5956
rect 6747 6012 6811 6016
rect 6747 5956 6751 6012
rect 6751 5956 6807 6012
rect 6807 5956 6811 6012
rect 6747 5952 6811 5956
rect 6827 6012 6891 6016
rect 6827 5956 6831 6012
rect 6831 5956 6887 6012
rect 6887 5956 6891 6012
rect 6827 5952 6891 5956
rect 6907 6012 6971 6016
rect 6907 5956 6911 6012
rect 6911 5956 6967 6012
rect 6967 5956 6971 6012
rect 6907 5952 6971 5956
rect 2428 5468 2492 5472
rect 2428 5412 2432 5468
rect 2432 5412 2488 5468
rect 2488 5412 2492 5468
rect 2428 5408 2492 5412
rect 2508 5468 2572 5472
rect 2508 5412 2512 5468
rect 2512 5412 2568 5468
rect 2568 5412 2572 5468
rect 2508 5408 2572 5412
rect 2588 5468 2652 5472
rect 2588 5412 2592 5468
rect 2592 5412 2648 5468
rect 2648 5412 2652 5468
rect 2588 5408 2652 5412
rect 2668 5468 2732 5472
rect 2668 5412 2672 5468
rect 2672 5412 2728 5468
rect 2728 5412 2732 5468
rect 2668 5408 2732 5412
rect 4061 5468 4125 5472
rect 4061 5412 4065 5468
rect 4065 5412 4121 5468
rect 4121 5412 4125 5468
rect 4061 5408 4125 5412
rect 4141 5468 4205 5472
rect 4141 5412 4145 5468
rect 4145 5412 4201 5468
rect 4201 5412 4205 5468
rect 4141 5408 4205 5412
rect 4221 5468 4285 5472
rect 4221 5412 4225 5468
rect 4225 5412 4281 5468
rect 4281 5412 4285 5468
rect 4221 5408 4285 5412
rect 4301 5468 4365 5472
rect 4301 5412 4305 5468
rect 4305 5412 4361 5468
rect 4361 5412 4365 5468
rect 4301 5408 4365 5412
rect 5694 5468 5758 5472
rect 5694 5412 5698 5468
rect 5698 5412 5754 5468
rect 5754 5412 5758 5468
rect 5694 5408 5758 5412
rect 5774 5468 5838 5472
rect 5774 5412 5778 5468
rect 5778 5412 5834 5468
rect 5834 5412 5838 5468
rect 5774 5408 5838 5412
rect 5854 5468 5918 5472
rect 5854 5412 5858 5468
rect 5858 5412 5914 5468
rect 5914 5412 5918 5468
rect 5854 5408 5918 5412
rect 5934 5468 5998 5472
rect 5934 5412 5938 5468
rect 5938 5412 5994 5468
rect 5994 5412 5998 5468
rect 5934 5408 5998 5412
rect 7327 5468 7391 5472
rect 7327 5412 7331 5468
rect 7331 5412 7387 5468
rect 7387 5412 7391 5468
rect 7327 5408 7391 5412
rect 7407 5468 7471 5472
rect 7407 5412 7411 5468
rect 7411 5412 7467 5468
rect 7467 5412 7471 5468
rect 7407 5408 7471 5412
rect 7487 5468 7551 5472
rect 7487 5412 7491 5468
rect 7491 5412 7547 5468
rect 7547 5412 7551 5468
rect 7487 5408 7551 5412
rect 7567 5468 7631 5472
rect 7567 5412 7571 5468
rect 7571 5412 7627 5468
rect 7627 5412 7631 5468
rect 7567 5408 7631 5412
rect 1768 4924 1832 4928
rect 1768 4868 1772 4924
rect 1772 4868 1828 4924
rect 1828 4868 1832 4924
rect 1768 4864 1832 4868
rect 1848 4924 1912 4928
rect 1848 4868 1852 4924
rect 1852 4868 1908 4924
rect 1908 4868 1912 4924
rect 1848 4864 1912 4868
rect 1928 4924 1992 4928
rect 1928 4868 1932 4924
rect 1932 4868 1988 4924
rect 1988 4868 1992 4924
rect 1928 4864 1992 4868
rect 2008 4924 2072 4928
rect 2008 4868 2012 4924
rect 2012 4868 2068 4924
rect 2068 4868 2072 4924
rect 2008 4864 2072 4868
rect 3401 4924 3465 4928
rect 3401 4868 3405 4924
rect 3405 4868 3461 4924
rect 3461 4868 3465 4924
rect 3401 4864 3465 4868
rect 3481 4924 3545 4928
rect 3481 4868 3485 4924
rect 3485 4868 3541 4924
rect 3541 4868 3545 4924
rect 3481 4864 3545 4868
rect 3561 4924 3625 4928
rect 3561 4868 3565 4924
rect 3565 4868 3621 4924
rect 3621 4868 3625 4924
rect 3561 4864 3625 4868
rect 3641 4924 3705 4928
rect 3641 4868 3645 4924
rect 3645 4868 3701 4924
rect 3701 4868 3705 4924
rect 3641 4864 3705 4868
rect 5034 4924 5098 4928
rect 5034 4868 5038 4924
rect 5038 4868 5094 4924
rect 5094 4868 5098 4924
rect 5034 4864 5098 4868
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 6667 4924 6731 4928
rect 6667 4868 6671 4924
rect 6671 4868 6727 4924
rect 6727 4868 6731 4924
rect 6667 4864 6731 4868
rect 6747 4924 6811 4928
rect 6747 4868 6751 4924
rect 6751 4868 6807 4924
rect 6807 4868 6811 4924
rect 6747 4864 6811 4868
rect 6827 4924 6891 4928
rect 6827 4868 6831 4924
rect 6831 4868 6887 4924
rect 6887 4868 6891 4924
rect 6827 4864 6891 4868
rect 6907 4924 6971 4928
rect 6907 4868 6911 4924
rect 6911 4868 6967 4924
rect 6967 4868 6971 4924
rect 6907 4864 6971 4868
rect 2428 4380 2492 4384
rect 2428 4324 2432 4380
rect 2432 4324 2488 4380
rect 2488 4324 2492 4380
rect 2428 4320 2492 4324
rect 2508 4380 2572 4384
rect 2508 4324 2512 4380
rect 2512 4324 2568 4380
rect 2568 4324 2572 4380
rect 2508 4320 2572 4324
rect 2588 4380 2652 4384
rect 2588 4324 2592 4380
rect 2592 4324 2648 4380
rect 2648 4324 2652 4380
rect 2588 4320 2652 4324
rect 2668 4380 2732 4384
rect 2668 4324 2672 4380
rect 2672 4324 2728 4380
rect 2728 4324 2732 4380
rect 2668 4320 2732 4324
rect 4061 4380 4125 4384
rect 4061 4324 4065 4380
rect 4065 4324 4121 4380
rect 4121 4324 4125 4380
rect 4061 4320 4125 4324
rect 4141 4380 4205 4384
rect 4141 4324 4145 4380
rect 4145 4324 4201 4380
rect 4201 4324 4205 4380
rect 4141 4320 4205 4324
rect 4221 4380 4285 4384
rect 4221 4324 4225 4380
rect 4225 4324 4281 4380
rect 4281 4324 4285 4380
rect 4221 4320 4285 4324
rect 4301 4380 4365 4384
rect 4301 4324 4305 4380
rect 4305 4324 4361 4380
rect 4361 4324 4365 4380
rect 4301 4320 4365 4324
rect 5694 4380 5758 4384
rect 5694 4324 5698 4380
rect 5698 4324 5754 4380
rect 5754 4324 5758 4380
rect 5694 4320 5758 4324
rect 5774 4380 5838 4384
rect 5774 4324 5778 4380
rect 5778 4324 5834 4380
rect 5834 4324 5838 4380
rect 5774 4320 5838 4324
rect 5854 4380 5918 4384
rect 5854 4324 5858 4380
rect 5858 4324 5914 4380
rect 5914 4324 5918 4380
rect 5854 4320 5918 4324
rect 5934 4380 5998 4384
rect 5934 4324 5938 4380
rect 5938 4324 5994 4380
rect 5994 4324 5998 4380
rect 5934 4320 5998 4324
rect 7327 4380 7391 4384
rect 7327 4324 7331 4380
rect 7331 4324 7387 4380
rect 7387 4324 7391 4380
rect 7327 4320 7391 4324
rect 7407 4380 7471 4384
rect 7407 4324 7411 4380
rect 7411 4324 7467 4380
rect 7467 4324 7471 4380
rect 7407 4320 7471 4324
rect 7487 4380 7551 4384
rect 7487 4324 7491 4380
rect 7491 4324 7547 4380
rect 7547 4324 7551 4380
rect 7487 4320 7551 4324
rect 7567 4380 7631 4384
rect 7567 4324 7571 4380
rect 7571 4324 7627 4380
rect 7627 4324 7631 4380
rect 7567 4320 7631 4324
rect 1768 3836 1832 3840
rect 1768 3780 1772 3836
rect 1772 3780 1828 3836
rect 1828 3780 1832 3836
rect 1768 3776 1832 3780
rect 1848 3836 1912 3840
rect 1848 3780 1852 3836
rect 1852 3780 1908 3836
rect 1908 3780 1912 3836
rect 1848 3776 1912 3780
rect 1928 3836 1992 3840
rect 1928 3780 1932 3836
rect 1932 3780 1988 3836
rect 1988 3780 1992 3836
rect 1928 3776 1992 3780
rect 2008 3836 2072 3840
rect 2008 3780 2012 3836
rect 2012 3780 2068 3836
rect 2068 3780 2072 3836
rect 2008 3776 2072 3780
rect 3401 3836 3465 3840
rect 3401 3780 3405 3836
rect 3405 3780 3461 3836
rect 3461 3780 3465 3836
rect 3401 3776 3465 3780
rect 3481 3836 3545 3840
rect 3481 3780 3485 3836
rect 3485 3780 3541 3836
rect 3541 3780 3545 3836
rect 3481 3776 3545 3780
rect 3561 3836 3625 3840
rect 3561 3780 3565 3836
rect 3565 3780 3621 3836
rect 3621 3780 3625 3836
rect 3561 3776 3625 3780
rect 3641 3836 3705 3840
rect 3641 3780 3645 3836
rect 3645 3780 3701 3836
rect 3701 3780 3705 3836
rect 3641 3776 3705 3780
rect 5034 3836 5098 3840
rect 5034 3780 5038 3836
rect 5038 3780 5094 3836
rect 5094 3780 5098 3836
rect 5034 3776 5098 3780
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 6667 3836 6731 3840
rect 6667 3780 6671 3836
rect 6671 3780 6727 3836
rect 6727 3780 6731 3836
rect 6667 3776 6731 3780
rect 6747 3836 6811 3840
rect 6747 3780 6751 3836
rect 6751 3780 6807 3836
rect 6807 3780 6811 3836
rect 6747 3776 6811 3780
rect 6827 3836 6891 3840
rect 6827 3780 6831 3836
rect 6831 3780 6887 3836
rect 6887 3780 6891 3836
rect 6827 3776 6891 3780
rect 6907 3836 6971 3840
rect 6907 3780 6911 3836
rect 6911 3780 6967 3836
rect 6967 3780 6971 3836
rect 6907 3776 6971 3780
rect 2428 3292 2492 3296
rect 2428 3236 2432 3292
rect 2432 3236 2488 3292
rect 2488 3236 2492 3292
rect 2428 3232 2492 3236
rect 2508 3292 2572 3296
rect 2508 3236 2512 3292
rect 2512 3236 2568 3292
rect 2568 3236 2572 3292
rect 2508 3232 2572 3236
rect 2588 3292 2652 3296
rect 2588 3236 2592 3292
rect 2592 3236 2648 3292
rect 2648 3236 2652 3292
rect 2588 3232 2652 3236
rect 2668 3292 2732 3296
rect 2668 3236 2672 3292
rect 2672 3236 2728 3292
rect 2728 3236 2732 3292
rect 2668 3232 2732 3236
rect 4061 3292 4125 3296
rect 4061 3236 4065 3292
rect 4065 3236 4121 3292
rect 4121 3236 4125 3292
rect 4061 3232 4125 3236
rect 4141 3292 4205 3296
rect 4141 3236 4145 3292
rect 4145 3236 4201 3292
rect 4201 3236 4205 3292
rect 4141 3232 4205 3236
rect 4221 3292 4285 3296
rect 4221 3236 4225 3292
rect 4225 3236 4281 3292
rect 4281 3236 4285 3292
rect 4221 3232 4285 3236
rect 4301 3292 4365 3296
rect 4301 3236 4305 3292
rect 4305 3236 4361 3292
rect 4361 3236 4365 3292
rect 4301 3232 4365 3236
rect 5694 3292 5758 3296
rect 5694 3236 5698 3292
rect 5698 3236 5754 3292
rect 5754 3236 5758 3292
rect 5694 3232 5758 3236
rect 5774 3292 5838 3296
rect 5774 3236 5778 3292
rect 5778 3236 5834 3292
rect 5834 3236 5838 3292
rect 5774 3232 5838 3236
rect 5854 3292 5918 3296
rect 5854 3236 5858 3292
rect 5858 3236 5914 3292
rect 5914 3236 5918 3292
rect 5854 3232 5918 3236
rect 5934 3292 5998 3296
rect 5934 3236 5938 3292
rect 5938 3236 5994 3292
rect 5994 3236 5998 3292
rect 5934 3232 5998 3236
rect 7327 3292 7391 3296
rect 7327 3236 7331 3292
rect 7331 3236 7387 3292
rect 7387 3236 7391 3292
rect 7327 3232 7391 3236
rect 7407 3292 7471 3296
rect 7407 3236 7411 3292
rect 7411 3236 7467 3292
rect 7467 3236 7471 3292
rect 7407 3232 7471 3236
rect 7487 3292 7551 3296
rect 7487 3236 7491 3292
rect 7491 3236 7547 3292
rect 7547 3236 7551 3292
rect 7487 3232 7551 3236
rect 7567 3292 7631 3296
rect 7567 3236 7571 3292
rect 7571 3236 7627 3292
rect 7627 3236 7631 3292
rect 7567 3232 7631 3236
rect 1768 2748 1832 2752
rect 1768 2692 1772 2748
rect 1772 2692 1828 2748
rect 1828 2692 1832 2748
rect 1768 2688 1832 2692
rect 1848 2748 1912 2752
rect 1848 2692 1852 2748
rect 1852 2692 1908 2748
rect 1908 2692 1912 2748
rect 1848 2688 1912 2692
rect 1928 2748 1992 2752
rect 1928 2692 1932 2748
rect 1932 2692 1988 2748
rect 1988 2692 1992 2748
rect 1928 2688 1992 2692
rect 2008 2748 2072 2752
rect 2008 2692 2012 2748
rect 2012 2692 2068 2748
rect 2068 2692 2072 2748
rect 2008 2688 2072 2692
rect 3401 2748 3465 2752
rect 3401 2692 3405 2748
rect 3405 2692 3461 2748
rect 3461 2692 3465 2748
rect 3401 2688 3465 2692
rect 3481 2748 3545 2752
rect 3481 2692 3485 2748
rect 3485 2692 3541 2748
rect 3541 2692 3545 2748
rect 3481 2688 3545 2692
rect 3561 2748 3625 2752
rect 3561 2692 3565 2748
rect 3565 2692 3621 2748
rect 3621 2692 3625 2748
rect 3561 2688 3625 2692
rect 3641 2748 3705 2752
rect 3641 2692 3645 2748
rect 3645 2692 3701 2748
rect 3701 2692 3705 2748
rect 3641 2688 3705 2692
rect 5034 2748 5098 2752
rect 5034 2692 5038 2748
rect 5038 2692 5094 2748
rect 5094 2692 5098 2748
rect 5034 2688 5098 2692
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 6667 2748 6731 2752
rect 6667 2692 6671 2748
rect 6671 2692 6727 2748
rect 6727 2692 6731 2748
rect 6667 2688 6731 2692
rect 6747 2748 6811 2752
rect 6747 2692 6751 2748
rect 6751 2692 6807 2748
rect 6807 2692 6811 2748
rect 6747 2688 6811 2692
rect 6827 2748 6891 2752
rect 6827 2692 6831 2748
rect 6831 2692 6887 2748
rect 6887 2692 6891 2748
rect 6827 2688 6891 2692
rect 6907 2748 6971 2752
rect 6907 2692 6911 2748
rect 6911 2692 6967 2748
rect 6967 2692 6971 2748
rect 6907 2688 6971 2692
rect 2428 2204 2492 2208
rect 2428 2148 2432 2204
rect 2432 2148 2488 2204
rect 2488 2148 2492 2204
rect 2428 2144 2492 2148
rect 2508 2204 2572 2208
rect 2508 2148 2512 2204
rect 2512 2148 2568 2204
rect 2568 2148 2572 2204
rect 2508 2144 2572 2148
rect 2588 2204 2652 2208
rect 2588 2148 2592 2204
rect 2592 2148 2648 2204
rect 2648 2148 2652 2204
rect 2588 2144 2652 2148
rect 2668 2204 2732 2208
rect 2668 2148 2672 2204
rect 2672 2148 2728 2204
rect 2728 2148 2732 2204
rect 2668 2144 2732 2148
rect 4061 2204 4125 2208
rect 4061 2148 4065 2204
rect 4065 2148 4121 2204
rect 4121 2148 4125 2204
rect 4061 2144 4125 2148
rect 4141 2204 4205 2208
rect 4141 2148 4145 2204
rect 4145 2148 4201 2204
rect 4201 2148 4205 2204
rect 4141 2144 4205 2148
rect 4221 2204 4285 2208
rect 4221 2148 4225 2204
rect 4225 2148 4281 2204
rect 4281 2148 4285 2204
rect 4221 2144 4285 2148
rect 4301 2204 4365 2208
rect 4301 2148 4305 2204
rect 4305 2148 4361 2204
rect 4361 2148 4365 2204
rect 4301 2144 4365 2148
rect 5694 2204 5758 2208
rect 5694 2148 5698 2204
rect 5698 2148 5754 2204
rect 5754 2148 5758 2204
rect 5694 2144 5758 2148
rect 5774 2204 5838 2208
rect 5774 2148 5778 2204
rect 5778 2148 5834 2204
rect 5834 2148 5838 2204
rect 5774 2144 5838 2148
rect 5854 2204 5918 2208
rect 5854 2148 5858 2204
rect 5858 2148 5914 2204
rect 5914 2148 5918 2204
rect 5854 2144 5918 2148
rect 5934 2204 5998 2208
rect 5934 2148 5938 2204
rect 5938 2148 5994 2204
rect 5994 2148 5998 2204
rect 5934 2144 5998 2148
rect 7327 2204 7391 2208
rect 7327 2148 7331 2204
rect 7331 2148 7387 2204
rect 7387 2148 7391 2204
rect 7327 2144 7391 2148
rect 7407 2204 7471 2208
rect 7407 2148 7411 2204
rect 7411 2148 7467 2204
rect 7467 2148 7471 2204
rect 7407 2144 7471 2148
rect 7487 2204 7551 2208
rect 7487 2148 7491 2204
rect 7491 2148 7547 2204
rect 7547 2148 7551 2204
rect 7487 2144 7551 2148
rect 7567 2204 7631 2208
rect 7567 2148 7571 2204
rect 7571 2148 7627 2204
rect 7627 2148 7631 2204
rect 7567 2144 7631 2148
<< metal4 >>
rect 1760 8192 2080 8752
rect 1760 8128 1768 8192
rect 1832 8128 1848 8192
rect 1912 8128 1928 8192
rect 1992 8128 2008 8192
rect 2072 8128 2080 8192
rect 1760 8006 2080 8128
rect 1760 7770 1802 8006
rect 2038 7770 2080 8006
rect 1760 7104 2080 7770
rect 1760 7040 1768 7104
rect 1832 7040 1848 7104
rect 1912 7040 1928 7104
rect 1992 7040 2008 7104
rect 2072 7040 2080 7104
rect 1760 6374 2080 7040
rect 1760 6138 1802 6374
rect 2038 6138 2080 6374
rect 1760 6016 2080 6138
rect 1760 5952 1768 6016
rect 1832 5952 1848 6016
rect 1912 5952 1928 6016
rect 1992 5952 2008 6016
rect 2072 5952 2080 6016
rect 1760 4928 2080 5952
rect 1760 4864 1768 4928
rect 1832 4864 1848 4928
rect 1912 4864 1928 4928
rect 1992 4864 2008 4928
rect 2072 4864 2080 4928
rect 1760 4742 2080 4864
rect 1760 4506 1802 4742
rect 2038 4506 2080 4742
rect 1760 3840 2080 4506
rect 1760 3776 1768 3840
rect 1832 3776 1848 3840
rect 1912 3776 1928 3840
rect 1992 3776 2008 3840
rect 2072 3776 2080 3840
rect 1760 3110 2080 3776
rect 1760 2874 1802 3110
rect 2038 2874 2080 3110
rect 1760 2752 2080 2874
rect 1760 2688 1768 2752
rect 1832 2688 1848 2752
rect 1912 2688 1928 2752
rect 1992 2688 2008 2752
rect 2072 2688 2080 2752
rect 1760 2128 2080 2688
rect 2420 8736 2740 8752
rect 2420 8672 2428 8736
rect 2492 8672 2508 8736
rect 2572 8672 2588 8736
rect 2652 8672 2668 8736
rect 2732 8672 2740 8736
rect 2420 8666 2740 8672
rect 2420 8430 2462 8666
rect 2698 8430 2740 8666
rect 2420 7648 2740 8430
rect 2420 7584 2428 7648
rect 2492 7584 2508 7648
rect 2572 7584 2588 7648
rect 2652 7584 2668 7648
rect 2732 7584 2740 7648
rect 2420 7034 2740 7584
rect 2420 6798 2462 7034
rect 2698 6798 2740 7034
rect 2420 6560 2740 6798
rect 2420 6496 2428 6560
rect 2492 6496 2508 6560
rect 2572 6496 2588 6560
rect 2652 6496 2668 6560
rect 2732 6496 2740 6560
rect 2420 5472 2740 6496
rect 2420 5408 2428 5472
rect 2492 5408 2508 5472
rect 2572 5408 2588 5472
rect 2652 5408 2668 5472
rect 2732 5408 2740 5472
rect 2420 5402 2740 5408
rect 2420 5166 2462 5402
rect 2698 5166 2740 5402
rect 2420 4384 2740 5166
rect 2420 4320 2428 4384
rect 2492 4320 2508 4384
rect 2572 4320 2588 4384
rect 2652 4320 2668 4384
rect 2732 4320 2740 4384
rect 2420 3770 2740 4320
rect 2420 3534 2462 3770
rect 2698 3534 2740 3770
rect 2420 3296 2740 3534
rect 2420 3232 2428 3296
rect 2492 3232 2508 3296
rect 2572 3232 2588 3296
rect 2652 3232 2668 3296
rect 2732 3232 2740 3296
rect 2420 2208 2740 3232
rect 2420 2144 2428 2208
rect 2492 2144 2508 2208
rect 2572 2144 2588 2208
rect 2652 2144 2668 2208
rect 2732 2144 2740 2208
rect 2420 2128 2740 2144
rect 3393 8192 3713 8752
rect 3393 8128 3401 8192
rect 3465 8128 3481 8192
rect 3545 8128 3561 8192
rect 3625 8128 3641 8192
rect 3705 8128 3713 8192
rect 3393 8006 3713 8128
rect 3393 7770 3435 8006
rect 3671 7770 3713 8006
rect 3393 7104 3713 7770
rect 3393 7040 3401 7104
rect 3465 7040 3481 7104
rect 3545 7040 3561 7104
rect 3625 7040 3641 7104
rect 3705 7040 3713 7104
rect 3393 6374 3713 7040
rect 3393 6138 3435 6374
rect 3671 6138 3713 6374
rect 3393 6016 3713 6138
rect 3393 5952 3401 6016
rect 3465 5952 3481 6016
rect 3545 5952 3561 6016
rect 3625 5952 3641 6016
rect 3705 5952 3713 6016
rect 3393 4928 3713 5952
rect 3393 4864 3401 4928
rect 3465 4864 3481 4928
rect 3545 4864 3561 4928
rect 3625 4864 3641 4928
rect 3705 4864 3713 4928
rect 3393 4742 3713 4864
rect 3393 4506 3435 4742
rect 3671 4506 3713 4742
rect 3393 3840 3713 4506
rect 3393 3776 3401 3840
rect 3465 3776 3481 3840
rect 3545 3776 3561 3840
rect 3625 3776 3641 3840
rect 3705 3776 3713 3840
rect 3393 3110 3713 3776
rect 3393 2874 3435 3110
rect 3671 2874 3713 3110
rect 3393 2752 3713 2874
rect 3393 2688 3401 2752
rect 3465 2688 3481 2752
rect 3545 2688 3561 2752
rect 3625 2688 3641 2752
rect 3705 2688 3713 2752
rect 3393 2128 3713 2688
rect 4053 8736 4373 8752
rect 4053 8672 4061 8736
rect 4125 8672 4141 8736
rect 4205 8672 4221 8736
rect 4285 8672 4301 8736
rect 4365 8672 4373 8736
rect 4053 8666 4373 8672
rect 4053 8430 4095 8666
rect 4331 8430 4373 8666
rect 4053 7648 4373 8430
rect 4053 7584 4061 7648
rect 4125 7584 4141 7648
rect 4205 7584 4221 7648
rect 4285 7584 4301 7648
rect 4365 7584 4373 7648
rect 4053 7034 4373 7584
rect 4053 6798 4095 7034
rect 4331 6798 4373 7034
rect 4053 6560 4373 6798
rect 4053 6496 4061 6560
rect 4125 6496 4141 6560
rect 4205 6496 4221 6560
rect 4285 6496 4301 6560
rect 4365 6496 4373 6560
rect 4053 5472 4373 6496
rect 4053 5408 4061 5472
rect 4125 5408 4141 5472
rect 4205 5408 4221 5472
rect 4285 5408 4301 5472
rect 4365 5408 4373 5472
rect 4053 5402 4373 5408
rect 4053 5166 4095 5402
rect 4331 5166 4373 5402
rect 4053 4384 4373 5166
rect 4053 4320 4061 4384
rect 4125 4320 4141 4384
rect 4205 4320 4221 4384
rect 4285 4320 4301 4384
rect 4365 4320 4373 4384
rect 4053 3770 4373 4320
rect 4053 3534 4095 3770
rect 4331 3534 4373 3770
rect 4053 3296 4373 3534
rect 4053 3232 4061 3296
rect 4125 3232 4141 3296
rect 4205 3232 4221 3296
rect 4285 3232 4301 3296
rect 4365 3232 4373 3296
rect 4053 2208 4373 3232
rect 4053 2144 4061 2208
rect 4125 2144 4141 2208
rect 4205 2144 4221 2208
rect 4285 2144 4301 2208
rect 4365 2144 4373 2208
rect 4053 2128 4373 2144
rect 5026 8192 5346 8752
rect 5026 8128 5034 8192
rect 5098 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5346 8192
rect 5026 8006 5346 8128
rect 5026 7770 5068 8006
rect 5304 7770 5346 8006
rect 5026 7104 5346 7770
rect 5026 7040 5034 7104
rect 5098 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5346 7104
rect 5026 6374 5346 7040
rect 5026 6138 5068 6374
rect 5304 6138 5346 6374
rect 5026 6016 5346 6138
rect 5026 5952 5034 6016
rect 5098 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5346 6016
rect 5026 4928 5346 5952
rect 5026 4864 5034 4928
rect 5098 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5346 4928
rect 5026 4742 5346 4864
rect 5026 4506 5068 4742
rect 5304 4506 5346 4742
rect 5026 3840 5346 4506
rect 5026 3776 5034 3840
rect 5098 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5346 3840
rect 5026 3110 5346 3776
rect 5026 2874 5068 3110
rect 5304 2874 5346 3110
rect 5026 2752 5346 2874
rect 5026 2688 5034 2752
rect 5098 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5346 2752
rect 5026 2128 5346 2688
rect 5686 8736 6006 8752
rect 5686 8672 5694 8736
rect 5758 8672 5774 8736
rect 5838 8672 5854 8736
rect 5918 8672 5934 8736
rect 5998 8672 6006 8736
rect 5686 8666 6006 8672
rect 5686 8430 5728 8666
rect 5964 8430 6006 8666
rect 5686 7648 6006 8430
rect 5686 7584 5694 7648
rect 5758 7584 5774 7648
rect 5838 7584 5854 7648
rect 5918 7584 5934 7648
rect 5998 7584 6006 7648
rect 5686 7034 6006 7584
rect 5686 6798 5728 7034
rect 5964 6798 6006 7034
rect 5686 6560 6006 6798
rect 5686 6496 5694 6560
rect 5758 6496 5774 6560
rect 5838 6496 5854 6560
rect 5918 6496 5934 6560
rect 5998 6496 6006 6560
rect 5686 5472 6006 6496
rect 5686 5408 5694 5472
rect 5758 5408 5774 5472
rect 5838 5408 5854 5472
rect 5918 5408 5934 5472
rect 5998 5408 6006 5472
rect 5686 5402 6006 5408
rect 5686 5166 5728 5402
rect 5964 5166 6006 5402
rect 5686 4384 6006 5166
rect 5686 4320 5694 4384
rect 5758 4320 5774 4384
rect 5838 4320 5854 4384
rect 5918 4320 5934 4384
rect 5998 4320 6006 4384
rect 5686 3770 6006 4320
rect 5686 3534 5728 3770
rect 5964 3534 6006 3770
rect 5686 3296 6006 3534
rect 5686 3232 5694 3296
rect 5758 3232 5774 3296
rect 5838 3232 5854 3296
rect 5918 3232 5934 3296
rect 5998 3232 6006 3296
rect 5686 2208 6006 3232
rect 5686 2144 5694 2208
rect 5758 2144 5774 2208
rect 5838 2144 5854 2208
rect 5918 2144 5934 2208
rect 5998 2144 6006 2208
rect 5686 2128 6006 2144
rect 6659 8192 6979 8752
rect 6659 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6907 8192
rect 6971 8128 6979 8192
rect 6659 8006 6979 8128
rect 6659 7770 6701 8006
rect 6937 7770 6979 8006
rect 6659 7104 6979 7770
rect 6659 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6907 7104
rect 6971 7040 6979 7104
rect 6659 6374 6979 7040
rect 6659 6138 6701 6374
rect 6937 6138 6979 6374
rect 6659 6016 6979 6138
rect 6659 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6907 6016
rect 6971 5952 6979 6016
rect 6659 4928 6979 5952
rect 6659 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6907 4928
rect 6971 4864 6979 4928
rect 6659 4742 6979 4864
rect 6659 4506 6701 4742
rect 6937 4506 6979 4742
rect 6659 3840 6979 4506
rect 6659 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6907 3840
rect 6971 3776 6979 3840
rect 6659 3110 6979 3776
rect 6659 2874 6701 3110
rect 6937 2874 6979 3110
rect 6659 2752 6979 2874
rect 6659 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6907 2752
rect 6971 2688 6979 2752
rect 6659 2128 6979 2688
rect 7319 8736 7639 8752
rect 7319 8672 7327 8736
rect 7391 8672 7407 8736
rect 7471 8672 7487 8736
rect 7551 8672 7567 8736
rect 7631 8672 7639 8736
rect 7319 8666 7639 8672
rect 7319 8430 7361 8666
rect 7597 8430 7639 8666
rect 7319 7648 7639 8430
rect 7319 7584 7327 7648
rect 7391 7584 7407 7648
rect 7471 7584 7487 7648
rect 7551 7584 7567 7648
rect 7631 7584 7639 7648
rect 7319 7034 7639 7584
rect 7319 6798 7361 7034
rect 7597 6798 7639 7034
rect 7319 6560 7639 6798
rect 7319 6496 7327 6560
rect 7391 6496 7407 6560
rect 7471 6496 7487 6560
rect 7551 6496 7567 6560
rect 7631 6496 7639 6560
rect 7319 5472 7639 6496
rect 7319 5408 7327 5472
rect 7391 5408 7407 5472
rect 7471 5408 7487 5472
rect 7551 5408 7567 5472
rect 7631 5408 7639 5472
rect 7319 5402 7639 5408
rect 7319 5166 7361 5402
rect 7597 5166 7639 5402
rect 7319 4384 7639 5166
rect 7319 4320 7327 4384
rect 7391 4320 7407 4384
rect 7471 4320 7487 4384
rect 7551 4320 7567 4384
rect 7631 4320 7639 4384
rect 7319 3770 7639 4320
rect 7319 3534 7361 3770
rect 7597 3534 7639 3770
rect 7319 3296 7639 3534
rect 7319 3232 7327 3296
rect 7391 3232 7407 3296
rect 7471 3232 7487 3296
rect 7551 3232 7567 3296
rect 7631 3232 7639 3296
rect 7319 2208 7639 3232
rect 7319 2144 7327 2208
rect 7391 2144 7407 2208
rect 7471 2144 7487 2208
rect 7551 2144 7567 2208
rect 7631 2144 7639 2208
rect 7319 2128 7639 2144
<< via4 >>
rect 1802 7770 2038 8006
rect 1802 6138 2038 6374
rect 1802 4506 2038 4742
rect 1802 2874 2038 3110
rect 2462 8430 2698 8666
rect 2462 6798 2698 7034
rect 2462 5166 2698 5402
rect 2462 3534 2698 3770
rect 3435 7770 3671 8006
rect 3435 6138 3671 6374
rect 3435 4506 3671 4742
rect 3435 2874 3671 3110
rect 4095 8430 4331 8666
rect 4095 6798 4331 7034
rect 4095 5166 4331 5402
rect 4095 3534 4331 3770
rect 5068 7770 5304 8006
rect 5068 6138 5304 6374
rect 5068 4506 5304 4742
rect 5068 2874 5304 3110
rect 5728 8430 5964 8666
rect 5728 6798 5964 7034
rect 5728 5166 5964 5402
rect 5728 3534 5964 3770
rect 6701 7770 6937 8006
rect 6701 6138 6937 6374
rect 6701 4506 6937 4742
rect 6701 2874 6937 3110
rect 7361 8430 7597 8666
rect 7361 6798 7597 7034
rect 7361 5166 7597 5402
rect 7361 3534 7597 3770
<< metal5 >>
rect 1056 8666 7684 8708
rect 1056 8430 2462 8666
rect 2698 8430 4095 8666
rect 4331 8430 5728 8666
rect 5964 8430 7361 8666
rect 7597 8430 7684 8666
rect 1056 8388 7684 8430
rect 1056 8006 7684 8048
rect 1056 7770 1802 8006
rect 2038 7770 3435 8006
rect 3671 7770 5068 8006
rect 5304 7770 6701 8006
rect 6937 7770 7684 8006
rect 1056 7728 7684 7770
rect 1056 7034 7684 7076
rect 1056 6798 2462 7034
rect 2698 6798 4095 7034
rect 4331 6798 5728 7034
rect 5964 6798 7361 7034
rect 7597 6798 7684 7034
rect 1056 6756 7684 6798
rect 1056 6374 7684 6416
rect 1056 6138 1802 6374
rect 2038 6138 3435 6374
rect 3671 6138 5068 6374
rect 5304 6138 6701 6374
rect 6937 6138 7684 6374
rect 1056 6096 7684 6138
rect 1056 5402 7684 5444
rect 1056 5166 2462 5402
rect 2698 5166 4095 5402
rect 4331 5166 5728 5402
rect 5964 5166 7361 5402
rect 7597 5166 7684 5402
rect 1056 5124 7684 5166
rect 1056 4742 7684 4784
rect 1056 4506 1802 4742
rect 2038 4506 3435 4742
rect 3671 4506 5068 4742
rect 5304 4506 6701 4742
rect 6937 4506 7684 4742
rect 1056 4464 7684 4506
rect 1056 3770 7684 3812
rect 1056 3534 2462 3770
rect 2698 3534 4095 3770
rect 4331 3534 5728 3770
rect 5964 3534 7361 3770
rect 7597 3534 7684 3770
rect 1056 3492 7684 3534
rect 1056 3110 7684 3152
rect 1056 2874 1802 3110
rect 2038 2874 3435 3110
rect 3671 2874 5068 3110
rect 5304 2874 6701 3110
rect 6937 2874 7684 3110
rect 1056 2832 7684 2874
use sky130_fd_sc_hd__inv_2  _30_
timestamp 0
transform -1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _31_
timestamp 0
transform -1 0 4968 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _32_
timestamp 0
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _33_
timestamp 0
transform 1 0 5152 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _34_
timestamp 0
transform 1 0 5244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _35_
timestamp 0
transform -1 0 6532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _36_
timestamp 0
transform -1 0 5336 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _37_
timestamp 0
transform 1 0 5428 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _38_
timestamp 0
transform -1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _39_
timestamp 0
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _40_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _41_
timestamp 0
transform -1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _42_
timestamp 0
transform 1 0 5520 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _43_
timestamp 0
transform -1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _44_
timestamp 0
transform 1 0 4968 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _45_
timestamp 0
transform -1 0 6072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _46_
timestamp 0
transform 1 0 4784 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _47_
timestamp 0
transform -1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _48_
timestamp 0
transform -1 0 2852 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _49_
timestamp 0
transform 1 0 2024 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _50_
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _51_
timestamp 0
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _52_
timestamp 0
transform -1 0 3864 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _53_
timestamp 0
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _54_
timestamp 0
transform 1 0 2576 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _55_
timestamp 0
transform 1 0 2668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _56_
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _57_
timestamp 0
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _58_
timestamp 0
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _59_
timestamp 0
transform 1 0 3864 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _60_
timestamp 0
transform -1 0 3680 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _61_
timestamp 0
transform 1 0 2392 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _62_
timestamp 0
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _63_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_20
timestamp 0
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 0
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65
timestamp 0
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_24
timestamp 0
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_36
timestamp 0
transform 1 0 4416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_44
timestamp 0
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_38
timestamp 0
transform 1 0 4600 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_59
timestamp 0
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_63
timestamp 0
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_20
timestamp 0
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_32
timestamp 0
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_44
timestamp 0
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_48
timestamp 0
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_65
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_37
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_46
timestamp 0
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_33
timestamp 0
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_38
timestamp 0
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_42
timestamp 0
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_46
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_63
timestamp 0
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_11
timestamp 0
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 0
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_18
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_22
timestamp 0
transform 1 0 3128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_30
timestamp 0
transform 1 0 3864 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_36
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_62
timestamp 0
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 0
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_37
timestamp 0
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_63
timestamp 0
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_67
timestamp 0
transform 1 0 7268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_12
timestamp 0
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_20
timestamp 0
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 0
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_63
timestamp 0
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_57
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_29
timestamp 0
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_37
timestamp 0
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 0
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_65
timestamp 0
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform -1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 0
transform -1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 0
transform -1 0 7360 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform -1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 0
transform -1 0 7360 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform -1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 7636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_26
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_28
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_29
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_30
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_31
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_32
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_33
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_34
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_35
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_36
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_37
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 4371 8704 4371 8704 4 VGND
rlabel metal1 s 4370 8160 4370 8160 4 VPWR
rlabel metal2 s 7314 2907 7314 2907 4 A[0]
rlabel metal2 s 7314 6239 7314 6239 4 A[1]
rlabel metal3 s 1050 6868 1050 6868 4 A[2]
rlabel metal2 s 3266 1588 3266 1588 4 A[3]
rlabel metal2 s 7222 5015 7222 5015 4 B[0]
rlabel metal1 s 7544 7854 7544 7854 4 B[1]
rlabel metal3 s 0 6128 800 6248 4 B[2]
port 7 nsew
rlabel metal2 s 2622 823 2622 823 4 B[3]
rlabel metal1 s 7544 5678 7544 5678 4 SEL[0]
rlabel metal1 s 7544 4590 7544 4590 4 SEL[1]
rlabel metal2 s 7222 3417 7222 3417 4 Y[0]
rlabel metal2 s 7222 7021 7222 7021 4 Y[1]
rlabel metal2 s 4002 9401 4002 9401 4 Y[2]
rlabel metal2 s 3910 1520 3910 1520 4 Y[3]
rlabel metal1 s 5658 6290 5658 6290 4 _00_
rlabel metal1 s 5014 3502 5014 3502 4 _01_
rlabel metal2 s 5750 3740 5750 3740 4 _02_
rlabel metal2 s 5474 3196 5474 3196 4 _03_
rlabel metal1 s 5336 6630 5336 6630 4 _04_
rlabel metal1 s 5106 5134 5106 5134 4 _05_
rlabel metal2 s 6118 5780 6118 5780 4 _06_
rlabel metal1 s 6118 6086 6118 6086 4 _07_
rlabel metal1 s 6118 6426 6118 6426 4 _08_
rlabel metal1 s 6486 6902 6486 6902 4 _09_
rlabel metal1 s 5980 6970 5980 6970 4 _10_
rlabel metal1 s 6854 6800 6854 6800 4 _11_
rlabel metal1 s 5520 6766 5520 6766 4 _12_
rlabel metal1 s 5198 6426 5198 6426 4 _13_
rlabel metal1 s 2645 7378 2645 7378 4 _14_
rlabel metal1 s 4370 5338 4370 5338 4 _15_
rlabel metal2 s 2162 6358 2162 6358 4 _16_
rlabel metal2 s 2622 6970 2622 6970 4 _17_
rlabel metal1 s 3128 7378 3128 7378 4 _18_
rlabel metal2 s 4002 6970 4002 6970 4 _19_
rlabel metal2 s 3818 6596 3818 6596 4 _20_
rlabel metal2 s 2990 3638 2990 3638 4 _21_
rlabel metal1 s 3266 6664 3266 6664 4 _22_
rlabel metal1 s 2806 3536 2806 3536 4 _23_
rlabel metal2 s 2898 3230 2898 3230 4 _24_
rlabel metal1 s 3174 3502 3174 3502 4 _25_
rlabel metal1 s 3726 3570 3726 3570 4 _26_
rlabel metal1 s 2714 3604 2714 3604 4 _27_
rlabel metal1 s 4002 3468 4002 3468 4 _28_
rlabel metal1 s 3542 3162 3542 3162 4 _29_
rlabel metal1 s 5750 2924 5750 2924 4 net1
rlabel metal1 s 6118 4794 6118 4794 4 net10
rlabel metal1 s 6164 3162 6164 3162 4 net11
rlabel metal2 s 6026 7106 6026 7106 4 net12
rlabel metal2 s 4462 7650 4462 7650 4 net13
rlabel metal1 s 4416 2414 4416 2414 4 net14
rlabel metal1 s 6808 6222 6808 6222 4 net2
rlabel metal1 s 2254 6800 2254 6800 4 net3
rlabel metal1 s 3082 2618 3082 2618 4 net4
rlabel metal1 s 6532 5270 6532 5270 4 net5
rlabel metal2 s 5750 6970 5750 6970 4 net6
rlabel metal1 s 1610 6188 1610 6188 4 net7
rlabel metal1 s 2392 3026 2392 3026 4 net8
rlabel metal1 s 4232 6358 4232 6358 4 net9
flabel metal3 s 8019 2728 8819 2848 0 FreeSans 600 0 0 0 A[0]
port 1 nsew
flabel metal3 s 8019 6128 8819 6248 0 FreeSans 600 0 0 0 A[1]
port 2 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 A[2]
port 3 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 A[3]
port 4 nsew
flabel metal3 s 8019 4768 8819 4888 0 FreeSans 600 0 0 0 B[0]
port 5 nsew
flabel metal3 s 8019 7488 8819 7608 0 FreeSans 600 0 0 0 B[1]
port 6 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 B[2]
flabel metal2 s 2594 0 2650 800 0 FreeSans 280 90 0 0 B[3]
port 8 nsew
flabel metal3 s 8019 5448 8819 5568 0 FreeSans 600 0 0 0 SEL[0]
port 9 nsew
flabel metal3 s 8019 4088 8819 4208 0 FreeSans 600 0 0 0 SEL[1]
port 10 nsew
flabel metal5 s 1056 8388 7684 8708 0 FreeSans 3200 0 0 0 VGND
port 11 nsew
flabel metal5 s 1056 6756 7684 7076 0 FreeSans 3200 0 0 0 VGND
port 11 nsew
flabel metal5 s 1056 5124 7684 5444 0 FreeSans 3200 0 0 0 VGND
port 11 nsew
flabel metal5 s 1056 3492 7684 3812 0 FreeSans 3200 0 0 0 VGND
port 11 nsew
flabel metal4 s 7319 2128 7639 8752 0 FreeSans 2400 90 0 0 VGND
port 11 nsew
flabel metal4 s 5686 2128 6006 8752 0 FreeSans 2400 90 0 0 VGND
port 11 nsew
flabel metal4 s 4053 2128 4373 8752 0 FreeSans 2400 90 0 0 VGND
port 11 nsew
flabel metal4 s 2420 2128 2740 8752 0 FreeSans 2400 90 0 0 VGND
port 11 nsew
flabel metal5 s 1056 7728 7684 8048 0 FreeSans 3200 0 0 0 VPWR
port 12 nsew
flabel metal5 s 1056 6096 7684 6416 0 FreeSans 3200 0 0 0 VPWR
port 12 nsew
flabel metal5 s 1056 4464 7684 4784 0 FreeSans 3200 0 0 0 VPWR
port 12 nsew
flabel metal5 s 1056 2832 7684 3152 0 FreeSans 3200 0 0 0 VPWR
port 12 nsew
flabel metal4 s 6659 2128 6979 8752 0 FreeSans 2400 90 0 0 VPWR
port 12 nsew
flabel metal4 s 5026 2128 5346 8752 0 FreeSans 2400 90 0 0 VPWR
port 12 nsew
flabel metal4 s 3393 2128 3713 8752 0 FreeSans 2400 90 0 0 VPWR
port 12 nsew
flabel metal4 s 1760 2128 2080 8752 0 FreeSans 2400 90 0 0 VPWR
port 12 nsew
flabel metal3 s 8019 3408 8819 3528 0 FreeSans 600 0 0 0 Y[0]
port 13 nsew
flabel metal3 s 8019 6808 8819 6928 0 FreeSans 600 0 0 0 Y[1]
port 14 nsew
flabel metal2 s 3882 10163 3938 10963 0 FreeSans 280 90 0 0 Y[2]
port 15 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 Y[3]
port 16 nsew
<< properties >>
string FIXED_BBOX 0 0 8819 10963
<< end >>
