module alu (A,
    B,
    SEL,
    Y);
 input [3:0] A;
 input [3:0] B;
 input [1:0] SEL;
 output [3:0] Y;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;

 sky130_fd_sc_hd__inv_2 _30_ (.A(SEL[1]),
    .Y(_00_));
 sky130_fd_sc_hd__or2_2 _31_ (.A(_00_),
    .B(SEL[0]),
    .X(_01_));
 sky130_fd_sc_hd__nand2_2 _32_ (.A(A[0]),
    .B(B[0]),
    .Y(_02_));
 sky130_fd_sc_hd__mux2_2 _33_ (.A0(SEL[1]),
    .A1(_01_),
    .S(_02_),
    .X(_03_));
 sky130_fd_sc_hd__o21a_2 _34_ (.A1(A[0]),
    .A2(B[0]),
    .B1(_03_),
    .X(Y[0]));
 sky130_fd_sc_hd__or2b_2 _35_ (.A(A[0]),
    .B_N(B[0]),
    .X(_04_));
 sky130_fd_sc_hd__or2b_2 _36_ (.A(SEL[1]),
    .B_N(SEL[0]),
    .X(_05_));
 sky130_fd_sc_hd__and3_2 _37_ (.A(B[0]),
    .B(B[1]),
    .C(_05_),
    .X(_06_));
 sky130_fd_sc_hd__a21oi_2 _38_ (.A1(B[0]),
    .A2(_05_),
    .B1(B[1]),
    .Y(_07_));
 sky130_fd_sc_hd__o21a_2 _39_ (.A1(_06_),
    .A2(_07_),
    .B1(A[1]),
    .X(_08_));
 sky130_fd_sc_hd__or3_2 _40_ (.A(A[1]),
    .B(_06_),
    .C(_07_),
    .X(_09_));
 sky130_fd_sc_hd__and2b_2 _41_ (.A_N(_08_),
    .B(_09_),
    .X(_10_));
 sky130_fd_sc_hd__xnor2_2 _42_ (.A(_04_),
    .B(_10_),
    .Y(_11_));
 sky130_fd_sc_hd__nand2_2 _43_ (.A(_00_),
    .B(_11_),
    .Y(_12_));
 sky130_fd_sc_hd__a211o_2 _44_ (.A1(SEL[0]),
    .A2(B[1]),
    .B1(A[1]),
    .C1(_00_),
    .X(_13_));
 sky130_fd_sc_hd__o211a_2 _45_ (.A1(B[1]),
    .A2(_01_),
    .B1(_12_),
    .C1(_13_),
    .X(Y[1]));
 sky130_fd_sc_hd__a21o_2 _46_ (.A1(_04_),
    .A2(_09_),
    .B1(_08_),
    .X(_14_));
 sky130_fd_sc_hd__o21ai_2 _47_ (.A1(B[0]),
    .A2(B[1]),
    .B1(_05_),
    .Y(_15_));
 sky130_fd_sc_hd__xnor2_2 _48_ (.A(B[2]),
    .B(_15_),
    .Y(_16_));
 sky130_fd_sc_hd__xnor2_2 _49_ (.A(A[2]),
    .B(_16_),
    .Y(_17_));
 sky130_fd_sc_hd__xnor2_2 _50_ (.A(_14_),
    .B(_17_),
    .Y(_18_));
 sky130_fd_sc_hd__nand2_2 _51_ (.A(_00_),
    .B(_18_),
    .Y(_19_));
 sky130_fd_sc_hd__a211o_2 _52_ (.A1(SEL[0]),
    .A2(A[2]),
    .B1(B[2]),
    .C1(_00_),
    .X(_20_));
 sky130_fd_sc_hd__o211a_2 _53_ (.A1(A[2]),
    .A2(_01_),
    .B1(_19_),
    .C1(_20_),
    .X(Y[2]));
 sky130_fd_sc_hd__and2_2 _54_ (.A(B[3]),
    .B(A[3]),
    .X(_21_));
 sky130_fd_sc_hd__and2b_2 _55_ (.A_N(_16_),
    .B(A[2]),
    .X(_22_));
 sky130_fd_sc_hd__a21oi_2 _56_ (.A1(_14_),
    .A2(_17_),
    .B1(_22_),
    .Y(_23_));
 sky130_fd_sc_hd__nor2_2 _57_ (.A(B[3]),
    .B(A[3]),
    .Y(_24_));
 sky130_fd_sc_hd__nor2_2 _58_ (.A(_24_),
    .B(_21_),
    .Y(_25_));
 sky130_fd_sc_hd__o31a_2 _59_ (.A1(B[0]),
    .A2(B[1]),
    .A3(B[2]),
    .B1(_05_),
    .X(_26_));
 sky130_fd_sc_hd__xnor2_2 _60_ (.A(_25_),
    .B(_26_),
    .Y(_27_));
 sky130_fd_sc_hd__xnor2_2 _61_ (.A(_23_),
    .B(_27_),
    .Y(_28_));
 sky130_fd_sc_hd__nand2_2 _62_ (.A(SEL[1]),
    .B(_24_),
    .Y(_29_));
 sky130_fd_sc_hd__o221a_2 _63_ (.A1(_01_),
    .A2(_21_),
    .B1(_28_),
    .B2(SEL[1]),
    .C1(_29_),
    .X(Y[3]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_37 ();
endmodule
