magic
tech sky130A
magscale 1 2
timestamp 1752153285
<< nwell >>
rect 1066 2159 7674 8721
<< obsli1 >>
rect 1104 2159 7636 8721
<< obsm1 >>
rect 842 2128 7806 8752
<< metal2 >>
rect 3882 10163 3938 10963
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
<< obsm2 >>
rect 846 10107 3826 10282
rect 3994 10107 7802 10282
rect 846 856 7802 10107
rect 846 734 2538 856
rect 2706 734 3182 856
rect 3350 734 3826 856
rect 3994 734 7802 856
<< metal3 >>
rect 8019 7488 8819 7608
rect 0 6808 800 6928
rect 8019 6808 8819 6928
rect 0 6128 800 6248
rect 8019 6128 8819 6248
rect 8019 5448 8819 5568
rect 8019 4768 8819 4888
rect 8019 4088 8819 4208
rect 8019 3408 8819 3528
rect 8019 2728 8819 2848
<< obsm3 >>
rect 798 7688 8019 8737
rect 798 7408 7939 7688
rect 798 7008 8019 7408
rect 880 6728 7939 7008
rect 798 6328 8019 6728
rect 880 6048 7939 6328
rect 798 5648 8019 6048
rect 798 5368 7939 5648
rect 798 4968 8019 5368
rect 798 4688 7939 4968
rect 798 4288 8019 4688
rect 798 4008 7939 4288
rect 798 3608 8019 4008
rect 798 3328 7939 3608
rect 798 2928 8019 3328
rect 798 2648 7939 2928
rect 798 2143 8019 2648
<< metal4 >>
rect 1760 2128 2080 8752
rect 2420 2128 2740 8752
rect 3393 2128 3713 8752
rect 4053 2128 4373 8752
rect 5026 2128 5346 8752
rect 5686 2128 6006 8752
rect 6659 2128 6979 8752
rect 7319 2128 7639 8752
<< metal5 >>
rect 1056 8388 7684 8708
rect 1056 7728 7684 8048
rect 1056 6756 7684 7076
rect 1056 6096 7684 6416
rect 1056 5124 7684 5444
rect 1056 4464 7684 4784
rect 1056 3492 7684 3812
rect 1056 2832 7684 3152
<< labels >>
rlabel metal3 s 8019 2728 8819 2848 6 A[0]
port 1 nsew signal input
rlabel metal3 s 8019 6128 8819 6248 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 A[2]
port 3 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 A[3]
port 4 nsew signal input
rlabel metal3 s 8019 4768 8819 4888 6 B[0]
port 5 nsew signal input
rlabel metal3 s 8019 7488 8819 7608 6 B[1]
port 6 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 B[2]
port 7 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 B[3]
port 8 nsew signal input
rlabel metal3 s 8019 5448 8819 5568 6 SEL[0]
port 9 nsew signal input
rlabel metal3 s 8019 4088 8819 4208 6 SEL[1]
port 10 nsew signal input
rlabel metal4 s 2420 2128 2740 8752 6 VGND
port 11 nsew ground bidirectional
rlabel metal4 s 4053 2128 4373 8752 6 VGND
port 11 nsew ground bidirectional
rlabel metal4 s 5686 2128 6006 8752 6 VGND
port 11 nsew ground bidirectional
rlabel metal4 s 7319 2128 7639 8752 6 VGND
port 11 nsew ground bidirectional
rlabel metal5 s 1056 3492 7684 3812 6 VGND
port 11 nsew ground bidirectional
rlabel metal5 s 1056 5124 7684 5444 6 VGND
port 11 nsew ground bidirectional
rlabel metal5 s 1056 6756 7684 7076 6 VGND
port 11 nsew ground bidirectional
rlabel metal5 s 1056 8388 7684 8708 6 VGND
port 11 nsew ground bidirectional
rlabel metal4 s 1760 2128 2080 8752 6 VPWR
port 12 nsew power bidirectional
rlabel metal4 s 3393 2128 3713 8752 6 VPWR
port 12 nsew power bidirectional
rlabel metal4 s 5026 2128 5346 8752 6 VPWR
port 12 nsew power bidirectional
rlabel metal4 s 6659 2128 6979 8752 6 VPWR
port 12 nsew power bidirectional
rlabel metal5 s 1056 2832 7684 3152 6 VPWR
port 12 nsew power bidirectional
rlabel metal5 s 1056 4464 7684 4784 6 VPWR
port 12 nsew power bidirectional
rlabel metal5 s 1056 6096 7684 6416 6 VPWR
port 12 nsew power bidirectional
rlabel metal5 s 1056 7728 7684 8048 6 VPWR
port 12 nsew power bidirectional
rlabel metal3 s 8019 3408 8819 3528 6 Y[0]
port 13 nsew signal output
rlabel metal3 s 8019 6808 8819 6928 6 Y[1]
port 14 nsew signal output
rlabel metal2 s 3882 10163 3938 10963 6 Y[2]
port 15 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 Y[3]
port 16 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8819 10963
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 312220
string GDS_FILE /openlane/designs/alu/runs/RUN_2025.07.10_13.13.56/results/signoff/alu.magic.gds
string GDS_START 154156
<< end >>

